magic
tech sky130A
timestamp 1745991594
<< error_s >>
rect 14518 23867 14519 23889
rect 14561 23867 14562 23889
rect 14518 23866 14562 23867
rect 16076 23867 16077 23889
rect 16119 23867 16120 23889
rect 16076 23866 16120 23867
rect 20504 23867 20505 23889
rect 20547 23867 20548 23889
rect 20504 23866 20548 23867
rect 22882 23867 22883 23889
rect 22925 23867 22926 23889
rect 22882 23866 22926 23867
rect 23948 23867 23949 23889
rect 23991 23867 23992 23889
rect 23948 23866 23992 23867
rect 25178 23867 25179 23889
rect 25221 23867 25222 23889
rect 25178 23866 25222 23867
rect 31164 23867 31165 23889
rect 31207 23867 31208 23889
rect 31164 23866 31208 23867
rect 12714 23375 12715 23397
rect 12757 23375 12758 23397
rect 12714 23374 12758 23375
rect 14531 23356 14569 23367
rect 31691 23356 31729 23367
rect 12078 23355 12764 23356
rect 12781 23355 13997 23356
rect 14441 23338 14458 23356
rect 14534 23338 14551 23356
rect 14605 23338 14622 23356
rect 14701 23338 14718 23356
rect 14794 23338 14811 23356
rect 14865 23338 14882 23356
rect 14961 23338 14978 23356
rect 15054 23338 15071 23356
rect 15125 23338 15142 23356
rect 15221 23338 15238 23356
rect 15314 23338 15331 23356
rect 15385 23338 15402 23356
rect 15481 23338 15498 23356
rect 15574 23338 15591 23356
rect 15645 23338 15662 23356
rect 15741 23338 15758 23356
rect 15834 23338 15851 23356
rect 15905 23338 15922 23356
rect 16001 23338 16018 23356
rect 16094 23338 16111 23356
rect 16165 23338 16182 23356
rect 16261 23338 16278 23356
rect 16354 23338 16371 23356
rect 16425 23338 16442 23356
rect 16521 23338 16538 23356
rect 16614 23338 16631 23356
rect 16685 23338 16702 23356
rect 16781 23338 16798 23356
rect 16874 23338 16891 23356
rect 16945 23338 16962 23356
rect 17041 23338 17058 23356
rect 17134 23338 17151 23356
rect 17205 23338 17222 23356
rect 17301 23338 17318 23356
rect 17394 23338 17411 23356
rect 17465 23338 17482 23356
rect 17561 23338 17578 23356
rect 17654 23338 17671 23356
rect 17725 23338 17742 23356
rect 17821 23338 17838 23356
rect 17914 23338 17931 23356
rect 17985 23338 18002 23356
rect 18081 23338 18098 23356
rect 18174 23338 18191 23356
rect 18245 23338 18262 23356
rect 18341 23338 18358 23356
rect 18434 23338 18451 23356
rect 18505 23338 18522 23356
rect 18601 23338 18618 23356
rect 18694 23338 18711 23356
rect 18765 23338 18782 23356
rect 18861 23338 18878 23356
rect 18954 23338 18971 23356
rect 19025 23338 19042 23356
rect 19121 23338 19138 23356
rect 19214 23338 19231 23356
rect 19285 23338 19302 23356
rect 19381 23338 19398 23356
rect 19474 23338 19491 23356
rect 19545 23338 19562 23356
rect 19641 23338 19658 23356
rect 19734 23338 19751 23356
rect 19805 23338 19822 23356
rect 19901 23338 19918 23356
rect 19994 23338 20011 23356
rect 20065 23338 20082 23356
rect 20161 23338 20178 23356
rect 20254 23338 20271 23356
rect 20325 23338 20342 23356
rect 20421 23338 20438 23356
rect 20514 23338 20531 23356
rect 20585 23338 20602 23356
rect 20681 23338 20698 23356
rect 20774 23338 20791 23356
rect 20845 23338 20862 23356
rect 20941 23338 20958 23356
rect 21034 23338 21051 23356
rect 21105 23338 21122 23356
rect 21201 23338 21218 23356
rect 21294 23338 21311 23356
rect 21365 23338 21382 23356
rect 21461 23338 21478 23356
rect 21554 23338 21571 23356
rect 21625 23338 21642 23356
rect 21721 23338 21738 23356
rect 21814 23338 21831 23356
rect 21885 23338 21902 23356
rect 21981 23338 21998 23356
rect 22074 23338 22091 23356
rect 22145 23338 22162 23356
rect 22241 23338 22258 23356
rect 22334 23338 22351 23356
rect 22405 23338 22422 23356
rect 22501 23338 22518 23356
rect 22594 23338 22611 23356
rect 22665 23338 22682 23356
rect 22761 23338 22778 23356
rect 22854 23338 22871 23356
rect 22925 23338 22942 23356
rect 23021 23338 23038 23356
rect 23114 23338 23131 23356
rect 23185 23338 23202 23356
rect 23281 23338 23298 23356
rect 23374 23338 23391 23356
rect 23445 23338 23462 23356
rect 23541 23338 23558 23356
rect 23634 23338 23651 23356
rect 23705 23338 23722 23356
rect 23801 23338 23818 23356
rect 23894 23338 23911 23356
rect 23965 23338 23982 23356
rect 24061 23338 24078 23356
rect 24154 23338 24171 23356
rect 24225 23338 24242 23356
rect 24321 23338 24338 23356
rect 24414 23338 24431 23356
rect 24485 23338 24502 23356
rect 24581 23338 24598 23356
rect 24674 23338 24691 23356
rect 24745 23338 24762 23356
rect 24841 23338 24858 23356
rect 24934 23338 24951 23356
rect 25005 23338 25022 23356
rect 25101 23338 25118 23356
rect 25194 23338 25211 23356
rect 25265 23338 25282 23356
rect 25361 23338 25378 23356
rect 25454 23338 25471 23356
rect 25525 23338 25542 23356
rect 25621 23338 25638 23356
rect 25714 23338 25731 23356
rect 25785 23338 25802 23356
rect 25881 23338 25898 23356
rect 25974 23338 25991 23356
rect 26045 23338 26062 23356
rect 26141 23338 26158 23356
rect 26234 23338 26251 23356
rect 26305 23338 26322 23356
rect 26401 23338 26418 23356
rect 26494 23338 26511 23356
rect 26565 23338 26582 23356
rect 26661 23338 26678 23356
rect 26754 23338 26771 23356
rect 26825 23338 26842 23356
rect 26921 23338 26938 23356
rect 27014 23338 27031 23356
rect 27085 23338 27102 23356
rect 27181 23338 27198 23356
rect 27274 23338 27291 23356
rect 27345 23338 27362 23356
rect 27441 23338 27458 23356
rect 27534 23338 27551 23356
rect 27605 23338 27622 23356
rect 27701 23338 27718 23356
rect 27794 23338 27811 23356
rect 27865 23338 27882 23356
rect 27961 23338 27978 23356
rect 28054 23338 28071 23356
rect 28125 23338 28142 23356
rect 28221 23338 28238 23356
rect 28314 23338 28331 23356
rect 28385 23338 28402 23356
rect 28481 23338 28498 23356
rect 28574 23338 28591 23356
rect 28645 23338 28662 23356
rect 28741 23338 28758 23356
rect 28834 23338 28851 23356
rect 28905 23338 28922 23356
rect 29001 23338 29018 23356
rect 29094 23338 29111 23356
rect 29165 23338 29182 23356
rect 29261 23338 29278 23356
rect 29354 23338 29371 23356
rect 29425 23338 29442 23356
rect 29521 23338 29538 23356
rect 29614 23338 29631 23356
rect 29685 23338 29702 23356
rect 29781 23338 29798 23356
rect 29874 23338 29891 23356
rect 29945 23338 29962 23356
rect 30041 23338 30058 23356
rect 30134 23338 30151 23356
rect 30205 23338 30222 23356
rect 30301 23338 30318 23356
rect 30394 23338 30411 23356
rect 30465 23338 30482 23356
rect 30561 23338 30578 23356
rect 30654 23338 30671 23356
rect 30725 23338 30742 23356
rect 30821 23338 30838 23356
rect 30914 23338 30931 23356
rect 30985 23338 31002 23356
rect 31081 23338 31098 23356
rect 31174 23338 31191 23356
rect 31245 23338 31262 23356
rect 31341 23338 31358 23356
rect 31434 23338 31451 23356
rect 31505 23338 31522 23356
rect 31601 23338 31618 23356
rect 31694 23338 31711 23356
rect 31765 23338 31782 23356
rect 12796 23335 12840 23336
rect 12796 23313 12797 23335
rect 12839 23313 12840 23335
rect 14531 23327 14569 23338
rect 31691 23327 31729 23338
rect 12586 23285 12603 23302
rect 12645 23285 12662 23302
rect 12213 23265 12230 23282
rect 12331 23265 12348 23282
rect 12907 23265 12924 23282
rect 13025 23265 13042 23282
rect 13280 23265 13297 23282
rect 13349 23265 13366 23282
rect 13427 23265 13444 23282
rect 13505 23265 13522 23282
rect 13583 23265 13600 23282
rect 13661 23265 13678 23282
rect 13739 23265 13756 23282
rect 13817 23265 13834 23282
rect 13885 23265 13902 23282
rect 13419 23256 13451 23257
rect 13575 23256 13607 23257
rect 13731 23256 13763 23257
rect 13816 23240 13817 23248
rect 13402 23239 13468 23240
rect 13558 23239 13624 23240
rect 13714 23239 13780 23240
rect 12302 23210 12303 23225
rect 12723 23204 12728 23221
rect 12996 23210 12997 23225
rect 13856 23210 13857 23225
rect 12740 23187 12745 23204
rect 13591 23122 13600 23139
rect 13591 23121 13617 23122
rect 13871 23058 13872 23073
rect 13833 22995 13834 23003
rect 12317 22974 12318 22989
rect 13011 22974 13012 22989
rect 13366 22986 13391 22987
rect 13402 22986 13469 22987
rect 13480 22986 13505 22987
rect 13522 22986 13547 22987
rect 13558 22986 13625 22987
rect 13636 22986 13661 22987
rect 13678 22986 13703 22987
rect 13714 22986 13781 22987
rect 13792 22986 13817 22987
rect 12357 22969 12365 22970
rect 13051 22969 13059 22970
rect 13366 22969 13374 22970
rect 13419 22969 13452 22970
rect 13497 22969 13505 22970
rect 13522 22969 13530 22970
rect 13575 22969 13608 22970
rect 13653 22969 13661 22970
rect 13678 22969 13686 22970
rect 13731 22969 13764 22970
rect 13809 22969 13817 22970
rect 12364 22952 12374 22953
rect 12381 22935 12391 22953
rect 13058 22952 13068 22953
rect 13075 22935 13085 22953
rect 13280 22945 13297 22962
rect 13349 22945 13366 22962
rect 13427 22945 13444 22962
rect 13505 22945 13522 22962
rect 13583 22945 13600 22962
rect 13661 22945 13678 22962
rect 13739 22945 13756 22962
rect 13817 22945 13834 22962
rect 13885 22945 13902 22962
rect 12213 22903 12230 22920
rect 12272 22903 12289 22920
rect 12331 22903 12348 22920
rect 12586 22903 12603 22920
rect 12645 22903 12662 22920
rect 12907 22903 12924 22920
rect 12966 22903 12983 22920
rect 13025 22903 13042 22920
rect 14026 22883 14027 22905
rect 14069 22883 14070 22905
rect 14026 22882 14070 22883
rect 12244 22848 12259 22849
rect 12303 22848 12318 22849
rect 12617 22848 12632 22849
rect 12938 22848 12953 22849
rect 12997 22848 13012 22849
rect 13311 22848 13326 22849
rect 13389 22848 13404 22849
rect 13467 22848 13482 22849
rect 13545 22848 13560 22849
rect 13623 22848 13638 22849
rect 13701 22848 13716 22849
rect 13779 22848 13794 22849
rect 13857 22848 13872 22849
rect 12755 22846 12765 22847
rect 12772 22846 12782 22847
rect 12714 22843 12758 22844
rect 12714 22821 12715 22843
rect 12757 22821 12758 22843
rect 14456 22829 14473 22847
rect 14531 22817 14569 22859
rect 14581 22829 14598 22847
rect 14631 22829 14648 22847
rect 14716 22829 14733 22847
rect 14794 22829 14811 22847
rect 14841 22829 14858 22847
rect 14891 22829 14908 22847
rect 14976 22829 14993 22847
rect 15054 22829 15071 22847
rect 15101 22829 15118 22847
rect 15151 22829 15168 22847
rect 15236 22829 15253 22847
rect 15314 22829 15331 22847
rect 15361 22829 15378 22847
rect 15411 22829 15428 22847
rect 15496 22829 15513 22847
rect 15574 22829 15591 22847
rect 15621 22829 15638 22847
rect 15671 22829 15688 22847
rect 15756 22829 15773 22847
rect 15834 22829 15851 22847
rect 15881 22829 15898 22847
rect 15931 22829 15948 22847
rect 16016 22829 16033 22847
rect 16094 22829 16111 22847
rect 16141 22829 16158 22847
rect 16191 22829 16208 22847
rect 16276 22829 16293 22847
rect 16354 22829 16371 22847
rect 16401 22829 16418 22847
rect 16451 22829 16468 22847
rect 16536 22829 16553 22847
rect 16614 22829 16631 22847
rect 16661 22829 16678 22847
rect 16711 22829 16728 22847
rect 16796 22829 16813 22847
rect 16874 22829 16891 22847
rect 16921 22829 16938 22847
rect 16971 22829 16988 22847
rect 17056 22829 17073 22847
rect 17134 22829 17151 22847
rect 17181 22829 17198 22847
rect 17231 22829 17248 22847
rect 17316 22829 17333 22847
rect 17394 22829 17411 22847
rect 17441 22829 17458 22847
rect 17491 22829 17508 22847
rect 17576 22829 17593 22847
rect 17654 22829 17671 22847
rect 17701 22829 17718 22847
rect 17751 22829 17768 22847
rect 17836 22829 17853 22847
rect 17914 22829 17931 22847
rect 17961 22829 17978 22847
rect 18011 22829 18028 22847
rect 18096 22829 18113 22847
rect 18174 22829 18191 22847
rect 18221 22829 18238 22847
rect 18271 22829 18288 22847
rect 18356 22829 18373 22847
rect 18434 22829 18451 22847
rect 18481 22829 18498 22847
rect 18531 22829 18548 22847
rect 18616 22829 18633 22847
rect 18694 22829 18711 22847
rect 18741 22829 18758 22847
rect 18791 22829 18808 22847
rect 18876 22829 18893 22847
rect 18954 22829 18971 22847
rect 19001 22829 19018 22847
rect 19051 22829 19068 22847
rect 19136 22829 19153 22847
rect 19214 22829 19231 22847
rect 19261 22829 19278 22847
rect 19311 22829 19328 22847
rect 19396 22829 19413 22847
rect 19474 22829 19491 22847
rect 19521 22829 19538 22847
rect 19571 22829 19588 22847
rect 19656 22829 19673 22847
rect 19734 22829 19751 22847
rect 19781 22829 19798 22847
rect 19831 22829 19848 22847
rect 19916 22829 19933 22847
rect 19994 22829 20011 22847
rect 20041 22829 20058 22847
rect 20091 22829 20108 22847
rect 20176 22829 20193 22847
rect 20254 22829 20271 22847
rect 20301 22829 20318 22847
rect 20351 22829 20368 22847
rect 20436 22829 20453 22847
rect 20514 22829 20531 22847
rect 20561 22829 20578 22847
rect 20611 22829 20628 22847
rect 20696 22829 20713 22847
rect 20774 22829 20791 22847
rect 20821 22829 20838 22847
rect 20871 22829 20888 22847
rect 20956 22829 20973 22847
rect 21034 22829 21051 22847
rect 21081 22829 21098 22847
rect 21131 22829 21148 22847
rect 21216 22829 21233 22847
rect 21294 22829 21311 22847
rect 21341 22829 21358 22847
rect 21391 22829 21408 22847
rect 21476 22829 21493 22847
rect 21554 22829 21571 22847
rect 21601 22829 21618 22847
rect 21651 22829 21668 22847
rect 21736 22829 21753 22847
rect 21814 22829 21831 22847
rect 21861 22829 21878 22847
rect 21911 22829 21928 22847
rect 21996 22829 22013 22847
rect 22074 22829 22091 22847
rect 22121 22829 22138 22847
rect 22171 22829 22188 22847
rect 22256 22829 22273 22847
rect 22334 22829 22351 22847
rect 22381 22829 22398 22847
rect 22431 22829 22448 22847
rect 22516 22829 22533 22847
rect 22594 22829 22611 22847
rect 22641 22829 22658 22847
rect 22691 22829 22708 22847
rect 22776 22829 22793 22847
rect 22854 22829 22871 22847
rect 22901 22829 22918 22847
rect 22951 22829 22968 22847
rect 23036 22829 23053 22847
rect 23114 22829 23131 22847
rect 23161 22829 23178 22847
rect 23211 22829 23228 22847
rect 23296 22829 23313 22847
rect 23374 22829 23391 22847
rect 23421 22829 23438 22847
rect 23471 22829 23488 22847
rect 23556 22829 23573 22847
rect 23634 22829 23651 22847
rect 23681 22829 23698 22847
rect 23731 22829 23748 22847
rect 23816 22829 23833 22847
rect 23894 22829 23911 22847
rect 23941 22829 23958 22847
rect 23991 22829 24008 22847
rect 24076 22829 24093 22847
rect 24154 22829 24171 22847
rect 24201 22829 24218 22847
rect 24251 22829 24268 22847
rect 24336 22829 24353 22847
rect 24414 22829 24431 22847
rect 24461 22829 24478 22847
rect 24511 22829 24528 22847
rect 24596 22829 24613 22847
rect 24674 22829 24691 22847
rect 24721 22829 24738 22847
rect 24771 22829 24788 22847
rect 24856 22829 24873 22847
rect 24934 22829 24951 22847
rect 24981 22829 24998 22847
rect 25031 22829 25048 22847
rect 25116 22829 25133 22847
rect 25194 22829 25211 22847
rect 25241 22829 25258 22847
rect 25291 22829 25308 22847
rect 25376 22829 25393 22847
rect 25454 22829 25471 22847
rect 25501 22829 25518 22847
rect 25551 22829 25568 22847
rect 25636 22829 25653 22847
rect 25714 22829 25731 22847
rect 25761 22829 25778 22847
rect 25811 22829 25828 22847
rect 25896 22829 25913 22847
rect 25974 22829 25991 22847
rect 26021 22829 26038 22847
rect 26071 22829 26088 22847
rect 26156 22829 26173 22847
rect 26234 22829 26251 22847
rect 26281 22829 26298 22847
rect 26331 22829 26348 22847
rect 26416 22829 26433 22847
rect 26494 22829 26511 22847
rect 26541 22829 26558 22847
rect 26591 22829 26608 22847
rect 26676 22829 26693 22847
rect 26754 22829 26771 22847
rect 26801 22829 26818 22847
rect 26851 22829 26868 22847
rect 26936 22829 26953 22847
rect 27014 22829 27031 22847
rect 27061 22829 27078 22847
rect 27111 22829 27128 22847
rect 27196 22829 27213 22847
rect 27274 22829 27291 22847
rect 27321 22829 27338 22847
rect 27371 22829 27388 22847
rect 27456 22829 27473 22847
rect 27534 22829 27551 22847
rect 27581 22829 27598 22847
rect 27631 22829 27648 22847
rect 27716 22829 27733 22847
rect 27794 22829 27811 22847
rect 27841 22829 27858 22847
rect 27891 22829 27908 22847
rect 27976 22829 27993 22847
rect 28054 22829 28071 22847
rect 28101 22829 28118 22847
rect 28151 22829 28168 22847
rect 28236 22829 28253 22847
rect 28314 22829 28331 22847
rect 28361 22829 28378 22847
rect 28411 22829 28428 22847
rect 28496 22829 28513 22847
rect 28574 22829 28591 22847
rect 28621 22829 28638 22847
rect 28671 22829 28688 22847
rect 28756 22829 28773 22847
rect 28834 22829 28851 22847
rect 28881 22829 28898 22847
rect 28931 22829 28948 22847
rect 29016 22829 29033 22847
rect 29094 22829 29111 22847
rect 29141 22829 29158 22847
rect 29191 22829 29208 22847
rect 29276 22829 29293 22847
rect 29354 22829 29371 22847
rect 29401 22829 29418 22847
rect 29451 22829 29468 22847
rect 29536 22829 29553 22847
rect 29614 22829 29631 22847
rect 29661 22829 29678 22847
rect 29711 22829 29728 22847
rect 29796 22829 29813 22847
rect 29874 22829 29891 22847
rect 29921 22829 29938 22847
rect 29971 22829 29988 22847
rect 30056 22829 30073 22847
rect 30134 22829 30151 22847
rect 30181 22829 30198 22847
rect 30231 22829 30248 22847
rect 30316 22829 30333 22847
rect 30394 22829 30411 22847
rect 30441 22829 30458 22847
rect 30491 22829 30508 22847
rect 30576 22829 30593 22847
rect 30654 22829 30671 22847
rect 30701 22829 30718 22847
rect 30751 22829 30768 22847
rect 30836 22829 30853 22847
rect 30914 22829 30931 22847
rect 30961 22829 30978 22847
rect 31011 22829 31028 22847
rect 31096 22829 31113 22847
rect 31174 22829 31191 22847
rect 31221 22829 31238 22847
rect 31271 22829 31288 22847
rect 31356 22829 31373 22847
rect 31434 22829 31451 22847
rect 31481 22829 31498 22847
rect 31531 22829 31548 22847
rect 31616 22829 31633 22847
rect 31691 22817 31729 22859
rect 31741 22829 31758 22847
rect 31791 22829 31808 22847
rect 12213 22756 12230 22773
rect 12272 22756 12289 22773
rect 12331 22756 12348 22773
rect 12586 22756 12603 22773
rect 12645 22756 12662 22773
rect 12907 22756 12924 22773
rect 12966 22756 12983 22773
rect 13025 22756 13042 22773
rect 12381 22724 12391 22741
rect 13075 22724 13085 22741
rect 12364 22723 12391 22724
rect 13058 22723 13085 22724
rect 12302 22702 12303 22717
rect 12996 22702 12997 22717
rect 13280 22714 13297 22731
rect 13349 22714 13366 22731
rect 13427 22714 13444 22731
rect 13505 22714 13522 22731
rect 13583 22714 13600 22731
rect 13661 22714 13678 22731
rect 13739 22714 13756 22731
rect 13817 22714 13834 22731
rect 13885 22714 13902 22731
rect 13366 22706 13374 22707
rect 13419 22706 13452 22707
rect 13497 22706 13505 22707
rect 13522 22706 13530 22707
rect 13575 22706 13608 22707
rect 13653 22706 13661 22707
rect 13678 22706 13686 22707
rect 13731 22706 13764 22707
rect 13809 22706 13817 22707
rect 13816 22690 13817 22698
rect 13366 22689 13391 22690
rect 13402 22689 13469 22690
rect 13480 22689 13505 22690
rect 13522 22689 13547 22690
rect 13558 22689 13625 22690
rect 13636 22689 13661 22690
rect 13678 22689 13703 22690
rect 13714 22689 13781 22690
rect 13792 22689 13817 22690
rect 13856 22618 13857 22633
rect 13591 22572 13600 22589
rect 13591 22571 13617 22572
rect 12317 22466 12318 22481
rect 12740 22473 12745 22489
rect 12723 22456 12728 22472
rect 13011 22466 13012 22481
rect 13871 22466 13872 22481
rect 13833 22445 13834 22453
rect 13402 22436 13468 22437
rect 13558 22436 13624 22437
rect 13714 22436 13780 22437
rect 13419 22419 13451 22420
rect 13575 22419 13607 22420
rect 13731 22419 13763 22420
rect 12213 22394 12230 22411
rect 12331 22394 12348 22411
rect 12907 22394 12924 22411
rect 13025 22394 13042 22411
rect 13280 22394 13297 22411
rect 13349 22394 13366 22411
rect 13427 22394 13444 22411
rect 13505 22394 13522 22411
rect 13583 22394 13600 22411
rect 13661 22394 13678 22411
rect 13739 22394 13756 22411
rect 13817 22394 13834 22411
rect 13885 22394 13902 22411
rect 12586 22374 12603 22391
rect 12645 22374 12662 22391
rect 14531 22338 14569 22349
rect 31691 22338 31729 22349
rect 12078 22337 12205 22338
rect 12238 22337 12381 22338
rect 12414 22337 12578 22338
rect 12611 22337 12695 22338
rect 12728 22337 12764 22338
rect 12781 22337 12899 22338
rect 12932 22337 13075 22338
rect 13108 22337 13272 22338
rect 13305 22337 13419 22338
rect 13451 22337 13575 22338
rect 13607 22337 13731 22338
rect 13763 22337 13877 22338
rect 13910 22337 13935 22338
rect 13968 22337 13997 22338
rect 14441 22320 14458 22338
rect 14518 22309 14519 22331
rect 14534 22320 14551 22338
rect 14561 22320 14562 22331
rect 14605 22320 14622 22338
rect 14701 22320 14718 22338
rect 14794 22320 14811 22338
rect 14865 22320 14882 22338
rect 14961 22320 14978 22338
rect 15054 22320 15071 22338
rect 15125 22320 15142 22338
rect 15221 22320 15238 22338
rect 15314 22320 15331 22338
rect 15385 22320 15402 22338
rect 15481 22320 15498 22338
rect 15574 22320 15591 22338
rect 15645 22320 15662 22338
rect 15741 22320 15758 22338
rect 15834 22320 15851 22338
rect 15905 22320 15922 22338
rect 16001 22320 16018 22338
rect 16094 22320 16111 22338
rect 16165 22320 16182 22338
rect 16261 22320 16278 22338
rect 16354 22320 16371 22338
rect 16425 22320 16442 22338
rect 16521 22320 16538 22338
rect 16614 22320 16631 22338
rect 16685 22320 16702 22338
rect 16781 22320 16798 22338
rect 16874 22320 16891 22338
rect 16945 22320 16962 22338
rect 17041 22320 17058 22338
rect 17134 22320 17151 22338
rect 17205 22320 17222 22338
rect 17301 22320 17318 22338
rect 17394 22320 17411 22338
rect 17465 22320 17482 22338
rect 17561 22320 17578 22338
rect 17654 22320 17671 22338
rect 17725 22320 17742 22338
rect 17821 22320 17838 22338
rect 17914 22320 17931 22338
rect 17985 22320 18002 22338
rect 18081 22320 18098 22338
rect 18174 22320 18191 22338
rect 18245 22320 18262 22338
rect 18341 22320 18358 22338
rect 18434 22320 18451 22338
rect 18505 22320 18522 22338
rect 18601 22320 18618 22338
rect 18694 22320 18711 22338
rect 18765 22320 18782 22338
rect 18861 22320 18878 22338
rect 18954 22320 18971 22338
rect 19025 22320 19042 22338
rect 19121 22320 19138 22338
rect 19214 22320 19231 22338
rect 19285 22320 19302 22338
rect 19381 22320 19398 22338
rect 19474 22320 19491 22338
rect 19545 22320 19562 22338
rect 19641 22320 19658 22338
rect 19734 22320 19751 22338
rect 19805 22320 19822 22338
rect 19901 22320 19918 22338
rect 19994 22320 20011 22338
rect 20065 22320 20082 22338
rect 30301 22320 30318 22338
rect 30394 22320 30411 22338
rect 30465 22320 30482 22338
rect 30561 22320 30578 22338
rect 30654 22320 30671 22338
rect 30725 22320 30742 22338
rect 30821 22320 30838 22338
rect 30914 22320 30931 22338
rect 30985 22320 31002 22338
rect 31081 22320 31098 22338
rect 31174 22320 31191 22338
rect 31245 22320 31262 22338
rect 31341 22320 31358 22338
rect 31434 22320 31451 22338
rect 31505 22320 31522 22338
rect 31601 22320 31618 22338
rect 31694 22320 31711 22338
rect 31765 22320 31782 22338
rect 14531 22309 14569 22320
rect 31691 22309 31729 22320
rect 14518 22308 14562 22309
rect 12586 22267 12603 22284
rect 12645 22267 12662 22284
rect 12796 22269 12840 22270
rect 12213 22247 12230 22264
rect 12331 22247 12348 22264
rect 12796 22247 12797 22269
rect 12839 22247 12840 22269
rect 12907 22247 12924 22264
rect 13025 22247 13042 22264
rect 13280 22247 13297 22264
rect 13349 22247 13366 22264
rect 13427 22247 13444 22264
rect 13505 22247 13522 22264
rect 13583 22247 13600 22264
rect 13661 22247 13678 22264
rect 13739 22247 13756 22264
rect 13817 22247 13834 22264
rect 13885 22247 13902 22264
rect 13419 22238 13451 22239
rect 13575 22238 13607 22239
rect 13731 22238 13763 22239
rect 13816 22222 13817 22230
rect 13402 22221 13468 22222
rect 13558 22221 13624 22222
rect 13714 22221 13780 22222
rect 12302 22192 12303 22207
rect 12723 22186 12728 22203
rect 12996 22192 12997 22207
rect 13856 22192 13857 22207
rect 12740 22169 12745 22186
rect 13591 22104 13600 22121
rect 13591 22103 13617 22104
rect 13871 22040 13872 22055
rect 13833 21977 13834 21985
rect 12317 21956 12318 21971
rect 13011 21956 13012 21971
rect 13366 21968 13391 21969
rect 13402 21968 13469 21969
rect 13480 21968 13505 21969
rect 13522 21968 13547 21969
rect 13558 21968 13625 21969
rect 13636 21968 13661 21969
rect 13678 21968 13703 21969
rect 13714 21968 13781 21969
rect 13792 21968 13817 21969
rect 12357 21951 12365 21952
rect 13051 21951 13059 21952
rect 13366 21951 13374 21952
rect 13419 21951 13452 21952
rect 13497 21951 13505 21952
rect 13522 21951 13530 21952
rect 13575 21951 13608 21952
rect 13653 21951 13661 21952
rect 13678 21951 13686 21952
rect 13731 21951 13764 21952
rect 13809 21951 13817 21952
rect 12364 21934 12374 21935
rect 12381 21917 12391 21935
rect 13058 21934 13068 21935
rect 13075 21917 13085 21935
rect 13280 21927 13297 21944
rect 13349 21927 13366 21944
rect 13427 21927 13444 21944
rect 13505 21927 13522 21944
rect 13583 21927 13600 21944
rect 13661 21927 13678 21944
rect 13739 21927 13756 21944
rect 13817 21927 13834 21944
rect 13885 21927 13902 21944
rect 12213 21885 12230 21902
rect 12272 21885 12289 21902
rect 12331 21885 12348 21902
rect 12586 21885 12603 21902
rect 12645 21885 12662 21902
rect 12907 21885 12924 21902
rect 12966 21885 12983 21902
rect 13025 21885 13042 21902
rect 12244 21830 12259 21831
rect 12303 21830 12318 21831
rect 12617 21830 12632 21831
rect 12938 21830 12953 21831
rect 12997 21830 13012 21831
rect 13311 21830 13326 21831
rect 13389 21830 13404 21831
rect 13467 21830 13482 21831
rect 13545 21830 13560 21831
rect 13623 21830 13638 21831
rect 13701 21830 13716 21831
rect 13779 21830 13794 21831
rect 13857 21830 13872 21831
rect 12755 21828 12765 21829
rect 12772 21828 12782 21829
rect 14456 21811 14473 21829
rect 14531 21799 14569 21841
rect 14581 21811 14598 21829
rect 14631 21811 14648 21829
rect 14716 21811 14733 21829
rect 14794 21811 14811 21829
rect 14841 21811 14858 21829
rect 14891 21811 14908 21829
rect 14976 21811 14993 21829
rect 15054 21811 15071 21829
rect 15101 21811 15118 21829
rect 15151 21811 15168 21829
rect 15236 21811 15253 21829
rect 15314 21811 15331 21829
rect 15361 21811 15378 21829
rect 15411 21811 15428 21829
rect 15496 21811 15513 21829
rect 15574 21811 15591 21829
rect 15621 21811 15638 21829
rect 15671 21811 15688 21829
rect 15756 21811 15773 21829
rect 15834 21811 15851 21829
rect 15881 21811 15898 21829
rect 15931 21811 15948 21829
rect 16016 21811 16033 21829
rect 16094 21811 16111 21829
rect 16141 21811 16158 21829
rect 16191 21811 16208 21829
rect 16276 21811 16293 21829
rect 16354 21811 16371 21829
rect 16401 21811 16418 21829
rect 16451 21811 16468 21829
rect 16536 21811 16553 21829
rect 16614 21811 16631 21829
rect 16661 21811 16678 21829
rect 16711 21811 16728 21829
rect 16796 21811 16813 21829
rect 16874 21811 16891 21829
rect 16921 21811 16938 21829
rect 16971 21811 16988 21829
rect 17056 21811 17073 21829
rect 17134 21811 17151 21829
rect 17181 21811 17198 21829
rect 17231 21811 17248 21829
rect 17316 21811 17333 21829
rect 17394 21811 17411 21829
rect 17441 21811 17458 21829
rect 17491 21811 17508 21829
rect 17576 21811 17593 21829
rect 17654 21811 17671 21829
rect 17701 21811 17718 21829
rect 17751 21811 17768 21829
rect 17836 21811 17853 21829
rect 17914 21811 17931 21829
rect 17961 21811 17978 21829
rect 18011 21811 18028 21829
rect 18096 21811 18113 21829
rect 18174 21811 18191 21829
rect 18221 21811 18238 21829
rect 18271 21811 18288 21829
rect 18356 21811 18373 21829
rect 18434 21811 18451 21829
rect 18481 21811 18498 21829
rect 18531 21811 18548 21829
rect 18616 21811 18633 21829
rect 18694 21811 18711 21829
rect 18741 21811 18758 21829
rect 18791 21811 18808 21829
rect 18876 21811 18893 21829
rect 18954 21811 18971 21829
rect 19001 21811 19018 21829
rect 19051 21811 19068 21829
rect 19136 21811 19153 21829
rect 19214 21811 19231 21829
rect 19261 21811 19278 21829
rect 19311 21811 19328 21829
rect 19396 21811 19413 21829
rect 19474 21811 19491 21829
rect 19521 21811 19538 21829
rect 19571 21811 19588 21829
rect 19656 21811 19673 21829
rect 19734 21811 19751 21829
rect 19781 21811 19798 21829
rect 19831 21811 19848 21829
rect 19916 21811 19933 21829
rect 19994 21811 20011 21829
rect 20041 21811 20058 21829
rect 20091 21811 20108 21829
rect 30240 21811 30248 21829
rect 30316 21811 30333 21829
rect 30394 21811 30411 21829
rect 30441 21811 30458 21829
rect 30491 21811 30508 21829
rect 30576 21811 30593 21829
rect 30654 21811 30671 21829
rect 30701 21811 30718 21829
rect 30751 21811 30768 21829
rect 30836 21811 30853 21829
rect 30914 21811 30931 21829
rect 30961 21811 30978 21829
rect 31011 21811 31028 21829
rect 31096 21811 31113 21829
rect 31174 21811 31191 21829
rect 31221 21811 31238 21829
rect 31271 21811 31288 21829
rect 31356 21811 31373 21829
rect 31434 21811 31451 21829
rect 31481 21811 31498 21829
rect 31531 21811 31548 21829
rect 31616 21811 31633 21829
rect 31691 21799 31729 21841
rect 31741 21811 31758 21829
rect 31791 21811 31808 21829
rect 12213 21738 12230 21755
rect 12272 21738 12289 21755
rect 12331 21738 12348 21755
rect 12586 21738 12603 21755
rect 12645 21738 12662 21755
rect 12907 21738 12924 21755
rect 12966 21738 12983 21755
rect 13025 21738 13042 21755
rect 12381 21706 12391 21723
rect 13075 21706 13085 21723
rect 12364 21705 12391 21706
rect 13058 21705 13085 21706
rect 12302 21684 12303 21699
rect 12996 21684 12997 21699
rect 13280 21696 13297 21713
rect 13349 21696 13366 21713
rect 13427 21696 13444 21713
rect 13505 21696 13522 21713
rect 13583 21696 13600 21713
rect 13661 21696 13678 21713
rect 13739 21696 13756 21713
rect 13817 21696 13834 21713
rect 13885 21696 13902 21713
rect 13366 21688 13374 21689
rect 13419 21688 13452 21689
rect 13497 21688 13505 21689
rect 13522 21688 13530 21689
rect 13575 21688 13608 21689
rect 13653 21688 13661 21689
rect 13678 21688 13686 21689
rect 13731 21688 13764 21689
rect 13809 21688 13817 21689
rect 13816 21672 13817 21680
rect 13366 21671 13391 21672
rect 13402 21671 13469 21672
rect 13480 21671 13505 21672
rect 13522 21671 13547 21672
rect 13558 21671 13625 21672
rect 13636 21671 13661 21672
rect 13678 21671 13703 21672
rect 13714 21671 13781 21672
rect 13792 21671 13817 21672
rect 13856 21600 13857 21615
rect 13591 21554 13600 21571
rect 13591 21553 13617 21554
rect 12317 21448 12318 21463
rect 12740 21455 12745 21471
rect 12723 21438 12728 21454
rect 13011 21448 13012 21463
rect 13871 21448 13872 21463
rect 13833 21427 13834 21435
rect 13402 21418 13468 21419
rect 13558 21418 13624 21419
rect 13714 21418 13780 21419
rect 13419 21401 13451 21402
rect 13575 21401 13607 21402
rect 13731 21401 13763 21402
rect 12213 21376 12230 21393
rect 12331 21376 12348 21393
rect 12907 21376 12924 21393
rect 13025 21376 13042 21393
rect 13280 21376 13297 21393
rect 13349 21376 13366 21393
rect 13427 21376 13444 21393
rect 13505 21376 13522 21393
rect 13583 21376 13600 21393
rect 13661 21376 13678 21393
rect 13739 21376 13756 21393
rect 13817 21376 13834 21393
rect 13885 21376 13902 21393
rect 12586 21356 12603 21373
rect 12645 21356 12662 21373
rect 14026 21325 14027 21347
rect 14069 21325 14070 21347
rect 14026 21324 14070 21325
rect 14531 21320 14569 21331
rect 31691 21320 31729 21331
rect 31738 21325 31739 21347
rect 31781 21325 31782 21347
rect 31738 21324 31782 21325
rect 12078 21319 12205 21320
rect 12238 21319 12381 21320
rect 12414 21319 12578 21320
rect 12611 21319 12695 21320
rect 12728 21319 12764 21320
rect 12781 21319 12899 21320
rect 12932 21319 13075 21320
rect 13108 21319 13272 21320
rect 13305 21319 13419 21320
rect 13451 21319 13575 21320
rect 13607 21319 13731 21320
rect 13763 21319 13877 21320
rect 13910 21319 13935 21320
rect 13968 21319 13997 21320
rect 14441 21302 14458 21320
rect 14534 21302 14551 21320
rect 14605 21302 14622 21320
rect 14701 21302 14718 21320
rect 14794 21302 14811 21320
rect 14865 21302 14882 21320
rect 14961 21302 14978 21320
rect 15054 21302 15071 21320
rect 15125 21302 15142 21320
rect 15221 21302 15238 21320
rect 15314 21302 15331 21320
rect 15385 21302 15402 21320
rect 15481 21302 15498 21320
rect 15574 21302 15591 21320
rect 15645 21302 15662 21320
rect 15741 21302 15758 21320
rect 15834 21302 15851 21320
rect 15905 21302 15922 21320
rect 16001 21302 16018 21320
rect 16094 21302 16111 21320
rect 16165 21302 16182 21320
rect 16261 21302 16278 21320
rect 16354 21302 16371 21320
rect 16425 21302 16442 21320
rect 16521 21302 16538 21320
rect 16614 21302 16631 21320
rect 16685 21302 16702 21320
rect 16781 21302 16798 21320
rect 16874 21302 16891 21320
rect 16945 21302 16962 21320
rect 17041 21302 17058 21320
rect 17134 21302 17151 21320
rect 17205 21302 17222 21320
rect 17301 21302 17318 21320
rect 17394 21302 17411 21320
rect 17465 21302 17482 21320
rect 17561 21302 17578 21320
rect 17654 21302 17671 21320
rect 17725 21302 17742 21320
rect 17821 21302 17838 21320
rect 17914 21302 17931 21320
rect 17985 21302 18002 21320
rect 18081 21302 18098 21320
rect 18174 21302 18191 21320
rect 18245 21302 18262 21320
rect 18341 21302 18358 21320
rect 18434 21302 18451 21320
rect 18505 21302 18522 21320
rect 18601 21302 18618 21320
rect 18694 21302 18711 21320
rect 18765 21302 18782 21320
rect 18861 21302 18878 21320
rect 18954 21302 18971 21320
rect 19025 21302 19042 21320
rect 19121 21302 19138 21320
rect 19214 21302 19231 21320
rect 19285 21302 19302 21320
rect 19381 21302 19398 21320
rect 19474 21302 19491 21320
rect 19545 21302 19562 21320
rect 19641 21302 19658 21320
rect 19734 21302 19751 21320
rect 19805 21302 19822 21320
rect 19901 21302 19918 21320
rect 19994 21302 20011 21320
rect 20065 21302 20082 21320
rect 30301 21302 30318 21320
rect 30394 21302 30411 21320
rect 30465 21302 30482 21320
rect 30561 21302 30578 21320
rect 30654 21302 30671 21320
rect 30725 21302 30742 21320
rect 30821 21302 30838 21320
rect 30914 21302 30931 21320
rect 30985 21302 31002 21320
rect 31081 21302 31098 21320
rect 31174 21302 31191 21320
rect 31245 21302 31262 21320
rect 31341 21302 31358 21320
rect 31434 21302 31451 21320
rect 31505 21302 31522 21320
rect 31601 21302 31618 21320
rect 31694 21302 31711 21320
rect 31765 21302 31782 21320
rect 14531 21291 14569 21302
rect 31691 21291 31729 21302
rect 13862 21285 13906 21286
rect 12586 21249 12603 21266
rect 12645 21249 12662 21266
rect 13862 21263 13863 21285
rect 13905 21263 13906 21285
rect 12213 21229 12230 21246
rect 12331 21229 12348 21246
rect 12907 21229 12924 21246
rect 13025 21229 13042 21246
rect 13280 21229 13297 21246
rect 13349 21229 13366 21246
rect 13427 21229 13444 21246
rect 13505 21229 13522 21246
rect 13583 21229 13600 21246
rect 13661 21229 13678 21246
rect 13739 21229 13756 21246
rect 13817 21229 13834 21246
rect 13885 21229 13902 21246
rect 13419 21220 13451 21221
rect 13575 21220 13607 21221
rect 13731 21220 13763 21221
rect 13816 21204 13817 21212
rect 13402 21203 13468 21204
rect 13558 21203 13624 21204
rect 13714 21203 13780 21204
rect 12302 21174 12303 21189
rect 12723 21168 12728 21185
rect 12996 21174 12997 21189
rect 13856 21174 13857 21189
rect 12740 21151 12745 21168
rect 13591 21086 13600 21103
rect 13591 21085 13617 21086
rect 13871 21022 13872 21037
rect 13833 20959 13834 20967
rect 12317 20938 12318 20953
rect 13011 20938 13012 20953
rect 13366 20950 13391 20951
rect 13402 20950 13469 20951
rect 13480 20950 13505 20951
rect 13522 20950 13547 20951
rect 13558 20950 13625 20951
rect 13636 20950 13661 20951
rect 13678 20950 13703 20951
rect 13714 20950 13781 20951
rect 13792 20950 13817 20951
rect 12357 20933 12365 20934
rect 13051 20933 13059 20934
rect 13366 20933 13374 20934
rect 13419 20933 13452 20934
rect 13497 20933 13505 20934
rect 13522 20933 13530 20934
rect 13575 20933 13608 20934
rect 13653 20933 13661 20934
rect 13678 20933 13686 20934
rect 13731 20933 13764 20934
rect 13809 20933 13817 20934
rect 12364 20916 12374 20917
rect 12381 20899 12391 20917
rect 13058 20916 13068 20917
rect 13075 20899 13085 20917
rect 13280 20909 13297 20926
rect 13349 20909 13366 20926
rect 13427 20909 13444 20926
rect 13505 20909 13522 20926
rect 13583 20909 13600 20926
rect 13661 20909 13678 20926
rect 13739 20909 13756 20926
rect 13817 20909 13834 20926
rect 13885 20909 13902 20926
rect 12213 20867 12230 20884
rect 12272 20867 12289 20884
rect 12331 20867 12348 20884
rect 12586 20867 12603 20884
rect 12645 20867 12662 20884
rect 12907 20867 12924 20884
rect 12966 20867 12983 20884
rect 13025 20867 13042 20884
rect 12714 20833 12715 20855
rect 12757 20833 12758 20855
rect 12714 20832 12758 20833
rect 13944 20833 13945 20855
rect 13987 20833 13988 20855
rect 13944 20832 13988 20833
rect 12244 20812 12259 20813
rect 12303 20812 12318 20813
rect 12617 20812 12632 20813
rect 12938 20812 12953 20813
rect 12997 20812 13012 20813
rect 13311 20812 13326 20813
rect 13389 20812 13404 20813
rect 13467 20812 13482 20813
rect 13545 20812 13560 20813
rect 13623 20812 13638 20813
rect 13701 20812 13716 20813
rect 13779 20812 13794 20813
rect 13857 20812 13872 20813
rect 12755 20810 12765 20811
rect 12772 20810 12782 20811
rect 12714 20793 12758 20794
rect 12714 20771 12715 20793
rect 12757 20771 12758 20793
rect 14026 20793 14070 20794
rect 14456 20793 14473 20811
rect 14026 20771 14027 20793
rect 14069 20771 14070 20793
rect 14531 20781 14569 20823
rect 14581 20793 14598 20811
rect 14631 20793 14648 20811
rect 14716 20793 14733 20811
rect 14794 20793 14811 20811
rect 14841 20793 14858 20811
rect 14891 20793 14908 20811
rect 14976 20793 14993 20811
rect 15054 20793 15071 20811
rect 15101 20793 15118 20811
rect 15151 20793 15168 20811
rect 15236 20793 15253 20811
rect 15314 20793 15331 20811
rect 15361 20793 15378 20811
rect 15411 20793 15428 20811
rect 15496 20793 15513 20811
rect 15574 20793 15591 20811
rect 15621 20793 15638 20811
rect 15671 20793 15688 20811
rect 15756 20793 15773 20811
rect 15834 20793 15851 20811
rect 15881 20793 15898 20811
rect 15931 20793 15948 20811
rect 16016 20793 16033 20811
rect 16094 20793 16111 20811
rect 16141 20793 16158 20811
rect 16191 20793 16208 20811
rect 16276 20793 16293 20811
rect 16354 20793 16371 20811
rect 16401 20793 16418 20811
rect 16451 20793 16468 20811
rect 16536 20793 16553 20811
rect 16614 20793 16631 20811
rect 16661 20793 16678 20811
rect 16711 20793 16728 20811
rect 16796 20793 16813 20811
rect 16874 20793 16891 20811
rect 16921 20793 16938 20811
rect 16971 20793 16988 20811
rect 17056 20793 17073 20811
rect 17134 20793 17151 20811
rect 17181 20793 17198 20811
rect 17231 20793 17248 20811
rect 17316 20793 17333 20811
rect 17394 20793 17411 20811
rect 17441 20793 17458 20811
rect 17491 20793 17508 20811
rect 17576 20793 17593 20811
rect 17654 20793 17671 20811
rect 17701 20793 17718 20811
rect 17751 20793 17768 20811
rect 17836 20793 17853 20811
rect 17914 20793 17931 20811
rect 17961 20793 17978 20811
rect 18011 20793 18028 20811
rect 18096 20793 18113 20811
rect 18174 20793 18191 20811
rect 18221 20793 18238 20811
rect 18271 20793 18288 20811
rect 18356 20793 18373 20811
rect 18434 20793 18451 20811
rect 18481 20793 18498 20811
rect 18531 20793 18548 20811
rect 18616 20793 18633 20811
rect 18694 20793 18711 20811
rect 18741 20793 18758 20811
rect 18791 20793 18808 20811
rect 18876 20793 18893 20811
rect 18954 20793 18971 20811
rect 19001 20793 19018 20811
rect 19051 20793 19068 20811
rect 19136 20793 19153 20811
rect 19214 20793 19231 20811
rect 19261 20793 19278 20811
rect 19311 20793 19328 20811
rect 19396 20793 19413 20811
rect 19474 20793 19491 20811
rect 19521 20793 19538 20811
rect 19571 20793 19588 20811
rect 19656 20793 19673 20811
rect 19734 20793 19751 20811
rect 19781 20793 19798 20811
rect 19831 20793 19848 20811
rect 19916 20793 19933 20811
rect 19994 20793 20011 20811
rect 20041 20793 20058 20811
rect 20091 20793 20108 20811
rect 30240 20793 30248 20811
rect 30316 20793 30333 20811
rect 30394 20793 30411 20811
rect 30441 20793 30458 20811
rect 30491 20793 30508 20811
rect 30576 20793 30593 20811
rect 30654 20793 30671 20811
rect 30701 20793 30718 20811
rect 30751 20793 30768 20811
rect 30836 20793 30853 20811
rect 30914 20793 30931 20811
rect 30961 20793 30978 20811
rect 31011 20793 31028 20811
rect 31096 20793 31113 20811
rect 31174 20793 31191 20811
rect 31221 20793 31238 20811
rect 31271 20793 31288 20811
rect 31356 20793 31373 20811
rect 31434 20793 31451 20811
rect 31481 20793 31498 20811
rect 31531 20793 31548 20811
rect 31616 20793 31633 20811
rect 31691 20781 31729 20823
rect 31741 20793 31758 20811
rect 31791 20793 31808 20811
rect 12213 20720 12230 20737
rect 12272 20720 12289 20737
rect 12331 20720 12348 20737
rect 12586 20720 12603 20737
rect 12645 20720 12662 20737
rect 12907 20720 12924 20737
rect 12966 20720 12983 20737
rect 13025 20720 13042 20737
rect 12381 20688 12391 20705
rect 13075 20688 13085 20705
rect 12364 20687 12391 20688
rect 13058 20687 13085 20688
rect 12302 20666 12303 20681
rect 12996 20666 12997 20681
rect 13280 20678 13297 20695
rect 13349 20678 13366 20695
rect 13427 20678 13444 20695
rect 13505 20678 13522 20695
rect 13583 20678 13600 20695
rect 13661 20678 13678 20695
rect 13739 20678 13756 20695
rect 13817 20678 13834 20695
rect 13885 20678 13902 20695
rect 13366 20670 13374 20671
rect 13419 20670 13452 20671
rect 13497 20670 13505 20671
rect 13522 20670 13530 20671
rect 13575 20670 13608 20671
rect 13653 20670 13661 20671
rect 13678 20670 13686 20671
rect 13731 20670 13764 20671
rect 13809 20670 13817 20671
rect 13816 20654 13817 20662
rect 13366 20653 13391 20654
rect 13402 20653 13469 20654
rect 13480 20653 13505 20654
rect 13522 20653 13547 20654
rect 13558 20653 13625 20654
rect 13636 20653 13661 20654
rect 13678 20653 13703 20654
rect 13714 20653 13781 20654
rect 13792 20653 13817 20654
rect 13856 20582 13857 20597
rect 13591 20536 13600 20553
rect 13591 20535 13617 20536
rect 12317 20430 12318 20445
rect 12740 20437 12745 20453
rect 12723 20420 12728 20436
rect 13011 20430 13012 20445
rect 13871 20430 13872 20445
rect 13833 20409 13834 20417
rect 13402 20400 13468 20401
rect 13558 20400 13624 20401
rect 13714 20400 13780 20401
rect 13419 20383 13451 20384
rect 13575 20383 13607 20384
rect 13731 20383 13763 20384
rect 12213 20358 12230 20375
rect 12331 20358 12348 20375
rect 12586 20338 12603 20355
rect 12645 20338 12662 20355
rect 12796 20341 12797 20363
rect 12839 20341 12840 20363
rect 12907 20358 12924 20375
rect 13025 20358 13042 20375
rect 13280 20358 13297 20375
rect 13349 20358 13366 20375
rect 13427 20358 13444 20375
rect 13505 20358 13522 20375
rect 13583 20358 13600 20375
rect 13661 20358 13678 20375
rect 13739 20358 13756 20375
rect 13817 20358 13834 20375
rect 13885 20358 13902 20375
rect 12796 20340 12840 20341
rect 14531 20302 14569 20313
rect 31691 20302 31729 20313
rect 12078 20301 12205 20302
rect 12238 20301 12381 20302
rect 12414 20301 12578 20302
rect 12611 20301 12695 20302
rect 12728 20301 12764 20302
rect 12781 20301 12899 20302
rect 12932 20301 13075 20302
rect 13108 20301 13272 20302
rect 13305 20301 13419 20302
rect 13451 20301 13575 20302
rect 13607 20301 13731 20302
rect 13763 20301 13877 20302
rect 13910 20301 13935 20302
rect 13944 20301 13997 20302
rect 13944 20279 13945 20301
rect 13987 20279 13988 20301
rect 14441 20284 14458 20302
rect 14534 20284 14551 20302
rect 14605 20284 14622 20302
rect 14701 20284 14718 20302
rect 14794 20284 14811 20302
rect 14865 20284 14882 20302
rect 14961 20284 14978 20302
rect 15054 20284 15071 20302
rect 15125 20284 15142 20302
rect 15221 20284 15238 20302
rect 15314 20284 15331 20302
rect 15385 20284 15402 20302
rect 15481 20284 15498 20302
rect 15574 20284 15591 20302
rect 15645 20284 15662 20302
rect 15741 20284 15758 20302
rect 15834 20284 15851 20302
rect 15905 20284 15922 20302
rect 16001 20284 16018 20302
rect 16094 20284 16111 20302
rect 16165 20284 16182 20302
rect 16261 20284 16278 20302
rect 16354 20284 16371 20302
rect 16425 20284 16442 20302
rect 16521 20284 16538 20302
rect 16614 20284 16631 20302
rect 16685 20284 16702 20302
rect 16781 20284 16798 20302
rect 16874 20284 16891 20302
rect 16945 20284 16962 20302
rect 17041 20284 17058 20302
rect 17134 20284 17151 20302
rect 17205 20284 17222 20302
rect 17301 20284 17318 20302
rect 17394 20284 17411 20302
rect 17465 20284 17482 20302
rect 17561 20284 17578 20302
rect 17654 20284 17671 20302
rect 17725 20284 17742 20302
rect 17821 20284 17838 20302
rect 17914 20284 17931 20302
rect 17985 20284 18002 20302
rect 18081 20284 18098 20302
rect 18174 20284 18191 20302
rect 18245 20284 18262 20302
rect 18341 20284 18358 20302
rect 18434 20284 18451 20302
rect 18505 20284 18522 20302
rect 18601 20284 18618 20302
rect 18694 20284 18711 20302
rect 18765 20284 18782 20302
rect 18861 20284 18878 20302
rect 18954 20284 18971 20302
rect 19025 20284 19042 20302
rect 19121 20284 19138 20302
rect 19214 20284 19231 20302
rect 19285 20284 19302 20302
rect 19381 20284 19398 20302
rect 19474 20284 19491 20302
rect 19545 20284 19562 20302
rect 19641 20284 19658 20302
rect 19734 20284 19751 20302
rect 19805 20284 19822 20302
rect 19901 20284 19918 20302
rect 19994 20284 20011 20302
rect 20065 20284 20082 20302
rect 30301 20284 30318 20302
rect 30394 20284 30411 20302
rect 30465 20284 30482 20302
rect 30561 20284 30578 20302
rect 30654 20284 30671 20302
rect 30725 20284 30742 20302
rect 30821 20284 30838 20302
rect 30914 20284 30931 20302
rect 30985 20284 31002 20302
rect 31081 20284 31098 20302
rect 31174 20284 31191 20302
rect 31245 20284 31262 20302
rect 31341 20284 31358 20302
rect 31434 20284 31451 20302
rect 31505 20284 31522 20302
rect 31601 20284 31618 20302
rect 31694 20284 31711 20302
rect 31765 20284 31782 20302
rect 14531 20273 14569 20284
rect 31691 20273 31729 20284
rect 12586 20231 12603 20248
rect 12645 20231 12662 20248
rect 12213 20211 12230 20228
rect 12331 20211 12348 20228
rect 12907 20211 12924 20228
rect 13025 20211 13042 20228
rect 13280 20211 13297 20228
rect 13349 20211 13366 20228
rect 13427 20211 13444 20228
rect 13505 20211 13522 20228
rect 13583 20211 13600 20228
rect 13661 20211 13678 20228
rect 13739 20211 13756 20228
rect 13817 20211 13834 20228
rect 13885 20211 13902 20228
rect 13419 20202 13451 20203
rect 13575 20202 13607 20203
rect 13731 20202 13763 20203
rect 13816 20186 13817 20194
rect 13402 20185 13468 20186
rect 13558 20185 13624 20186
rect 13714 20185 13780 20186
rect 12302 20156 12303 20171
rect 12723 20150 12728 20167
rect 12996 20156 12997 20171
rect 13856 20156 13857 20171
rect 12740 20133 12745 20150
rect 13591 20068 13600 20085
rect 13591 20067 13617 20068
rect 13871 20004 13872 20019
rect 13833 19941 13834 19949
rect 12317 19920 12318 19935
rect 13011 19920 13012 19935
rect 13366 19932 13391 19933
rect 13402 19932 13469 19933
rect 13480 19932 13505 19933
rect 13522 19932 13547 19933
rect 13558 19932 13625 19933
rect 13636 19932 13661 19933
rect 13678 19932 13703 19933
rect 13714 19932 13781 19933
rect 13792 19932 13817 19933
rect 12357 19915 12365 19916
rect 13051 19915 13059 19916
rect 13366 19915 13374 19916
rect 13419 19915 13452 19916
rect 13497 19915 13505 19916
rect 13522 19915 13530 19916
rect 13575 19915 13608 19916
rect 13653 19915 13661 19916
rect 13678 19915 13686 19916
rect 13731 19915 13764 19916
rect 13809 19915 13817 19916
rect 12364 19898 12374 19899
rect 12381 19881 12391 19899
rect 13058 19898 13068 19899
rect 13075 19881 13085 19899
rect 13280 19891 13297 19908
rect 13349 19891 13366 19908
rect 13427 19891 13444 19908
rect 13505 19891 13522 19908
rect 13583 19891 13600 19908
rect 13661 19891 13678 19908
rect 13739 19891 13756 19908
rect 13817 19891 13834 19908
rect 13885 19891 13902 19908
rect 12213 19849 12230 19866
rect 12272 19849 12289 19866
rect 12331 19849 12348 19866
rect 12586 19849 12603 19866
rect 12645 19849 12662 19866
rect 12907 19849 12924 19866
rect 12966 19849 12983 19866
rect 13025 19849 13042 19866
rect 12244 19794 12259 19795
rect 12303 19794 12318 19795
rect 12617 19794 12632 19795
rect 12938 19794 12953 19795
rect 12997 19794 13012 19795
rect 13311 19794 13326 19795
rect 13389 19794 13404 19795
rect 13467 19794 13482 19795
rect 13545 19794 13560 19795
rect 13623 19794 13638 19795
rect 13701 19794 13716 19795
rect 13779 19794 13794 19795
rect 13857 19794 13872 19795
rect 12755 19792 12765 19793
rect 12772 19792 12782 19793
rect 14456 19775 14473 19793
rect 14531 19763 14569 19805
rect 14581 19775 14598 19793
rect 14631 19775 14648 19793
rect 14716 19775 14733 19793
rect 14794 19775 14811 19793
rect 14841 19775 14858 19793
rect 14891 19775 14908 19793
rect 14976 19775 14993 19793
rect 15054 19775 15071 19793
rect 15101 19775 15118 19793
rect 15151 19775 15168 19793
rect 15236 19775 15253 19793
rect 31022 19775 31028 19793
rect 31096 19775 31113 19793
rect 31174 19775 31191 19793
rect 31221 19775 31238 19793
rect 31271 19775 31288 19793
rect 31356 19775 31373 19793
rect 31434 19775 31451 19793
rect 31481 19775 31498 19793
rect 31531 19775 31548 19793
rect 31616 19775 31633 19793
rect 31691 19763 31729 19805
rect 31741 19775 31758 19793
rect 31791 19775 31808 19793
rect 12714 19727 12758 19728
rect 12213 19702 12230 19719
rect 12272 19702 12289 19719
rect 12331 19702 12348 19719
rect 12586 19702 12603 19719
rect 12645 19702 12662 19719
rect 12714 19705 12715 19727
rect 12757 19705 12758 19727
rect 12907 19702 12924 19719
rect 12966 19702 12983 19719
rect 13025 19702 13042 19719
rect 12381 19670 12391 19687
rect 13075 19670 13085 19687
rect 12364 19669 12391 19670
rect 13058 19669 13085 19670
rect 12302 19648 12303 19663
rect 12996 19648 12997 19663
rect 13280 19660 13297 19677
rect 13349 19660 13366 19677
rect 13427 19660 13444 19677
rect 13505 19660 13522 19677
rect 13583 19660 13600 19677
rect 13661 19660 13678 19677
rect 13739 19660 13756 19677
rect 13817 19660 13834 19677
rect 13885 19660 13902 19677
rect 13366 19652 13374 19653
rect 13419 19652 13452 19653
rect 13497 19652 13505 19653
rect 13522 19652 13530 19653
rect 13575 19652 13608 19653
rect 13653 19652 13661 19653
rect 13678 19652 13686 19653
rect 13731 19652 13764 19653
rect 13809 19652 13817 19653
rect 13816 19636 13817 19644
rect 13366 19635 13391 19636
rect 13402 19635 13469 19636
rect 13480 19635 13505 19636
rect 13522 19635 13547 19636
rect 13558 19635 13625 19636
rect 13636 19635 13661 19636
rect 13678 19635 13703 19636
rect 13714 19635 13781 19636
rect 13792 19635 13817 19636
rect 13856 19564 13857 19579
rect 13591 19518 13600 19535
rect 13591 19517 13617 19518
rect 12317 19412 12318 19427
rect 12740 19419 12745 19435
rect 12723 19402 12728 19418
rect 13011 19412 13012 19427
rect 13871 19412 13872 19427
rect 13833 19391 13834 19399
rect 13402 19382 13468 19383
rect 13558 19382 13624 19383
rect 13714 19382 13780 19383
rect 13419 19365 13451 19366
rect 13575 19365 13607 19366
rect 13731 19365 13763 19366
rect 12213 19340 12230 19357
rect 12331 19340 12348 19357
rect 12907 19340 12924 19357
rect 13025 19340 13042 19357
rect 13280 19340 13297 19357
rect 13349 19340 13366 19357
rect 13427 19340 13444 19357
rect 13505 19340 13522 19357
rect 13583 19340 13600 19357
rect 13661 19340 13678 19357
rect 13739 19340 13756 19357
rect 13817 19340 13834 19357
rect 13885 19340 13902 19357
rect 12586 19320 12603 19337
rect 12645 19320 12662 19337
rect 12796 19284 12797 19297
rect 12839 19284 12840 19297
rect 14531 19284 14569 19295
rect 31691 19284 31729 19295
rect 12078 19283 12205 19284
rect 12238 19283 12381 19284
rect 12414 19283 12578 19284
rect 12611 19283 12695 19284
rect 12728 19283 12764 19284
rect 12781 19283 12899 19284
rect 12932 19283 13075 19284
rect 13108 19283 13272 19284
rect 13305 19283 13419 19284
rect 13451 19283 13575 19284
rect 13607 19283 13731 19284
rect 13763 19283 13877 19284
rect 13910 19283 13935 19284
rect 13968 19283 13997 19284
rect 12796 19275 12797 19283
rect 12839 19275 12840 19283
rect 12796 19274 12840 19275
rect 14441 19266 14458 19284
rect 14534 19266 14551 19284
rect 14605 19266 14622 19284
rect 14701 19266 14718 19284
rect 14794 19266 14811 19284
rect 14865 19266 14882 19284
rect 14961 19266 14978 19284
rect 15054 19266 15071 19284
rect 15125 19266 15142 19284
rect 15221 19266 15238 19284
rect 31081 19266 31098 19284
rect 31174 19266 31191 19284
rect 31245 19266 31262 19284
rect 31341 19266 31358 19284
rect 31434 19266 31451 19284
rect 31505 19266 31522 19284
rect 31601 19266 31618 19284
rect 31694 19266 31711 19284
rect 31765 19266 31782 19284
rect 14531 19255 14569 19266
rect 31691 19255 31729 19266
rect 12796 19235 12840 19236
rect 12586 19213 12603 19230
rect 12645 19213 12662 19230
rect 12796 19213 12797 19235
rect 12839 19213 12840 19235
rect 14518 19235 14562 19236
rect 14518 19213 14519 19235
rect 14561 19213 14562 19235
rect 31738 19235 31782 19236
rect 31738 19213 31739 19235
rect 31781 19213 31782 19235
rect 12213 19193 12230 19210
rect 12331 19193 12348 19210
rect 12907 19193 12924 19210
rect 13025 19193 13042 19210
rect 13280 19193 13297 19210
rect 13349 19193 13366 19210
rect 13427 19193 13444 19210
rect 13505 19193 13522 19210
rect 13583 19193 13600 19210
rect 13661 19193 13678 19210
rect 13739 19193 13756 19210
rect 13817 19193 13834 19210
rect 13885 19193 13902 19210
rect 13419 19184 13451 19185
rect 13575 19184 13607 19185
rect 13731 19184 13763 19185
rect 13816 19168 13817 19176
rect 13402 19167 13468 19168
rect 13558 19167 13624 19168
rect 13714 19167 13780 19168
rect 12302 19138 12303 19153
rect 12723 19132 12728 19149
rect 12996 19138 12997 19153
rect 13856 19138 13857 19153
rect 12740 19115 12745 19132
rect 13591 19050 13600 19067
rect 13591 19049 13617 19050
rect 13871 18986 13872 19001
rect 13833 18923 13834 18931
rect 12317 18902 12318 18917
rect 13011 18902 13012 18917
rect 13366 18914 13391 18915
rect 13402 18914 13469 18915
rect 13480 18914 13505 18915
rect 13522 18914 13547 18915
rect 13558 18914 13625 18915
rect 13636 18914 13661 18915
rect 13678 18914 13703 18915
rect 13714 18914 13781 18915
rect 13792 18914 13817 18915
rect 12357 18897 12365 18898
rect 13051 18897 13059 18898
rect 13366 18897 13374 18898
rect 13419 18897 13452 18898
rect 13497 18897 13505 18898
rect 13522 18897 13530 18898
rect 13575 18897 13608 18898
rect 13653 18897 13661 18898
rect 13678 18897 13686 18898
rect 13731 18897 13764 18898
rect 13809 18897 13817 18898
rect 12364 18880 12374 18881
rect 12381 18863 12391 18881
rect 13058 18880 13068 18881
rect 13075 18863 13085 18881
rect 13280 18873 13297 18890
rect 13349 18873 13366 18890
rect 13427 18873 13444 18890
rect 13505 18873 13522 18890
rect 13583 18873 13600 18890
rect 13661 18873 13678 18890
rect 13739 18873 13756 18890
rect 13817 18873 13834 18890
rect 13885 18873 13902 18890
rect 12213 18831 12230 18848
rect 12272 18831 12289 18848
rect 12331 18831 12348 18848
rect 12586 18831 12603 18848
rect 12645 18831 12662 18848
rect 12907 18831 12924 18848
rect 12966 18831 12983 18848
rect 13025 18831 13042 18848
rect 12244 18776 12259 18777
rect 12303 18776 12318 18777
rect 12617 18776 12632 18777
rect 12938 18776 12953 18777
rect 12997 18776 13012 18777
rect 13311 18776 13326 18777
rect 13389 18776 13404 18777
rect 13467 18776 13482 18777
rect 13545 18776 13560 18777
rect 13623 18776 13638 18777
rect 13701 18776 13716 18777
rect 13779 18776 13794 18777
rect 13857 18776 13872 18777
rect 12755 18774 12765 18775
rect 12772 18774 12782 18775
rect 14456 18757 14473 18775
rect 14531 18745 14569 18787
rect 14600 18783 14601 18805
rect 14643 18783 14644 18805
rect 14600 18782 14644 18783
rect 14581 18757 14598 18775
rect 14631 18757 14648 18775
rect 14716 18757 14733 18775
rect 14794 18757 14811 18775
rect 14841 18757 14858 18775
rect 14891 18757 14908 18775
rect 14976 18757 14993 18775
rect 15054 18757 15071 18775
rect 15101 18757 15118 18775
rect 15151 18757 15168 18775
rect 15236 18757 15253 18775
rect 31022 18757 31028 18775
rect 31096 18757 31113 18775
rect 31174 18757 31191 18775
rect 31221 18757 31238 18775
rect 31271 18757 31288 18775
rect 31356 18757 31373 18775
rect 31434 18757 31451 18775
rect 31481 18757 31498 18775
rect 31531 18757 31548 18775
rect 31616 18757 31633 18775
rect 31691 18745 31729 18787
rect 31741 18757 31758 18775
rect 31791 18757 31808 18775
rect 14026 18743 14070 18744
rect 14026 18721 14027 18743
rect 14069 18721 14070 18743
rect 12213 18684 12230 18701
rect 12272 18684 12289 18701
rect 12331 18684 12348 18701
rect 12586 18684 12603 18701
rect 12645 18684 12662 18701
rect 12907 18684 12924 18701
rect 12966 18684 12983 18701
rect 13025 18684 13042 18701
rect 12381 18652 12391 18669
rect 13075 18652 13085 18669
rect 12364 18651 12391 18652
rect 13058 18651 13085 18652
rect 12302 18630 12303 18645
rect 12996 18630 12997 18645
rect 13280 18642 13297 18659
rect 13349 18642 13366 18659
rect 13427 18642 13444 18659
rect 13505 18642 13522 18659
rect 13583 18642 13600 18659
rect 13661 18642 13678 18659
rect 13739 18642 13756 18659
rect 13817 18642 13834 18659
rect 13885 18642 13902 18659
rect 13366 18634 13374 18635
rect 13419 18634 13452 18635
rect 13497 18634 13505 18635
rect 13522 18634 13530 18635
rect 13575 18634 13608 18635
rect 13653 18634 13661 18635
rect 13678 18634 13686 18635
rect 13731 18634 13764 18635
rect 13809 18634 13817 18635
rect 13816 18618 13817 18626
rect 13366 18617 13391 18618
rect 13402 18617 13469 18618
rect 13480 18617 13505 18618
rect 13522 18617 13547 18618
rect 13558 18617 13625 18618
rect 13636 18617 13661 18618
rect 13678 18617 13703 18618
rect 13714 18617 13781 18618
rect 13792 18617 13817 18618
rect 13856 18546 13857 18561
rect 13591 18500 13600 18517
rect 13591 18499 13617 18500
rect 12317 18394 12318 18409
rect 12740 18401 12745 18417
rect 12723 18384 12728 18400
rect 13011 18394 13012 18409
rect 13871 18394 13872 18409
rect 13833 18373 13834 18381
rect 13402 18364 13468 18365
rect 13558 18364 13624 18365
rect 13714 18364 13780 18365
rect 13419 18347 13451 18348
rect 13575 18347 13607 18348
rect 13731 18347 13763 18348
rect 12213 18322 12230 18339
rect 12331 18322 12348 18339
rect 12907 18322 12924 18339
rect 13025 18322 13042 18339
rect 13280 18322 13297 18339
rect 13349 18322 13366 18339
rect 13427 18322 13444 18339
rect 13505 18322 13522 18339
rect 13583 18322 13600 18339
rect 13661 18322 13678 18339
rect 13739 18322 13756 18339
rect 13817 18322 13834 18339
rect 13885 18322 13902 18339
rect 12586 18302 12603 18319
rect 12645 18302 12662 18319
rect 14531 18266 14569 18277
rect 31691 18266 31729 18277
rect 12078 18265 12205 18266
rect 12238 18265 12381 18266
rect 12414 18265 12578 18266
rect 12611 18265 12695 18266
rect 12728 18265 12764 18266
rect 12781 18265 12899 18266
rect 12932 18265 13075 18266
rect 13108 18265 13272 18266
rect 13305 18265 13419 18266
rect 13451 18265 13575 18266
rect 13607 18265 13731 18266
rect 13763 18265 13877 18266
rect 13910 18265 13935 18266
rect 13968 18265 13997 18266
rect 14108 18251 14152 18252
rect 14108 18229 14109 18251
rect 14151 18229 14152 18251
rect 14441 18248 14458 18266
rect 14534 18248 14551 18266
rect 14605 18248 14622 18266
rect 14701 18248 14718 18266
rect 14794 18248 14811 18266
rect 14865 18248 14882 18266
rect 14961 18248 14978 18266
rect 15054 18248 15071 18266
rect 15125 18248 15142 18266
rect 15221 18248 15238 18266
rect 31081 18248 31098 18266
rect 31174 18248 31191 18266
rect 31245 18248 31262 18266
rect 31341 18248 31358 18266
rect 31434 18248 31451 18266
rect 31505 18248 31522 18266
rect 31601 18248 31618 18266
rect 31694 18248 31711 18266
rect 31765 18248 31782 18266
rect 14531 18237 14569 18248
rect 31691 18237 31729 18248
rect 12586 18195 12603 18212
rect 12645 18195 12662 18212
rect 12213 18175 12230 18192
rect 12331 18175 12348 18192
rect 12907 18175 12924 18192
rect 13025 18175 13042 18192
rect 13280 18175 13297 18192
rect 13349 18175 13366 18192
rect 13427 18175 13444 18192
rect 13505 18175 13522 18192
rect 13583 18175 13600 18192
rect 13661 18175 13678 18192
rect 13739 18175 13756 18192
rect 13817 18175 13834 18192
rect 13885 18175 13902 18192
rect 13419 18166 13451 18167
rect 13575 18166 13607 18167
rect 13731 18166 13763 18167
rect 13816 18150 13817 18158
rect 13402 18149 13468 18150
rect 13558 18149 13624 18150
rect 13714 18149 13780 18150
rect 12302 18120 12303 18135
rect 12723 18114 12728 18131
rect 12996 18120 12997 18135
rect 13856 18120 13857 18135
rect 12740 18097 12745 18114
rect 13591 18032 13600 18049
rect 13591 18031 13617 18032
rect 13871 17968 13872 17983
rect 13833 17905 13834 17913
rect 12317 17884 12318 17899
rect 13011 17884 13012 17899
rect 13366 17896 13391 17897
rect 13402 17896 13469 17897
rect 13480 17896 13505 17897
rect 13522 17896 13547 17897
rect 13558 17896 13625 17897
rect 13636 17896 13661 17897
rect 13678 17896 13703 17897
rect 13714 17896 13781 17897
rect 13792 17896 13817 17897
rect 12357 17879 12365 17880
rect 13051 17879 13059 17880
rect 13366 17879 13374 17880
rect 13419 17879 13452 17880
rect 13497 17879 13505 17880
rect 13522 17879 13530 17880
rect 13575 17879 13608 17880
rect 13653 17879 13661 17880
rect 13678 17879 13686 17880
rect 13731 17879 13764 17880
rect 13809 17879 13817 17880
rect 12364 17862 12374 17863
rect 12381 17845 12391 17863
rect 13058 17862 13068 17863
rect 13075 17845 13085 17863
rect 13280 17855 13297 17872
rect 13349 17855 13366 17872
rect 13427 17855 13444 17872
rect 13505 17855 13522 17872
rect 13583 17855 13600 17872
rect 13661 17855 13678 17872
rect 13739 17855 13756 17872
rect 13817 17855 13834 17872
rect 13885 17855 13902 17872
rect 12213 17813 12230 17830
rect 12272 17813 12289 17830
rect 12331 17813 12348 17830
rect 12586 17813 12603 17830
rect 12645 17813 12662 17830
rect 12714 17799 12715 17821
rect 12757 17799 12758 17821
rect 12907 17813 12924 17830
rect 12966 17813 12983 17830
rect 13025 17813 13042 17830
rect 12714 17798 12758 17799
rect 12714 17759 12758 17760
rect 13944 17759 13988 17760
rect 12244 17758 12259 17759
rect 12303 17758 12318 17759
rect 12617 17758 12632 17759
rect 12714 17737 12715 17759
rect 12757 17757 12758 17759
rect 12938 17758 12953 17759
rect 12997 17758 13012 17759
rect 13311 17758 13326 17759
rect 13389 17758 13404 17759
rect 13467 17758 13482 17759
rect 13545 17758 13560 17759
rect 13623 17758 13638 17759
rect 13701 17758 13716 17759
rect 13779 17758 13794 17759
rect 13857 17758 13872 17759
rect 12755 17756 12765 17757
rect 12772 17756 12782 17757
rect 12757 17737 12758 17756
rect 13944 17737 13945 17759
rect 13987 17737 13988 17759
rect 14456 17739 14473 17757
rect 14531 17727 14569 17769
rect 14581 17739 14598 17757
rect 14631 17739 14648 17757
rect 14716 17739 14733 17757
rect 14794 17739 14811 17757
rect 14841 17739 14858 17757
rect 14891 17739 14908 17757
rect 14976 17739 14993 17757
rect 15054 17739 15071 17757
rect 15101 17739 15118 17757
rect 15151 17739 15168 17757
rect 15236 17739 15253 17757
rect 31022 17739 31028 17757
rect 31096 17739 31113 17757
rect 31174 17739 31191 17757
rect 31221 17739 31238 17757
rect 31271 17739 31288 17757
rect 31356 17739 31373 17757
rect 31434 17739 31451 17757
rect 31481 17739 31498 17757
rect 31531 17739 31548 17757
rect 31616 17739 31633 17757
rect 31691 17727 31729 17769
rect 31741 17739 31758 17757
rect 31791 17739 31808 17757
rect 12213 17666 12230 17683
rect 12272 17666 12289 17683
rect 12331 17666 12348 17683
rect 12586 17666 12603 17683
rect 12645 17666 12662 17683
rect 12907 17666 12924 17683
rect 12966 17666 12983 17683
rect 13025 17666 13042 17683
rect 12381 17634 12391 17651
rect 13075 17634 13085 17651
rect 12364 17633 12391 17634
rect 13058 17633 13085 17634
rect 12302 17612 12303 17627
rect 12996 17612 12997 17627
rect 13280 17624 13297 17641
rect 13349 17624 13366 17641
rect 13427 17624 13444 17641
rect 13505 17624 13522 17641
rect 13583 17624 13600 17641
rect 13661 17624 13678 17641
rect 13739 17624 13756 17641
rect 13817 17624 13834 17641
rect 13885 17624 13902 17641
rect 13366 17616 13374 17617
rect 13419 17616 13452 17617
rect 13497 17616 13505 17617
rect 13522 17616 13530 17617
rect 13575 17616 13608 17617
rect 13653 17616 13661 17617
rect 13678 17616 13686 17617
rect 13731 17616 13764 17617
rect 13809 17616 13817 17617
rect 13816 17600 13817 17608
rect 13366 17599 13391 17600
rect 13402 17599 13469 17600
rect 13480 17599 13505 17600
rect 13522 17599 13547 17600
rect 13558 17599 13625 17600
rect 13636 17599 13661 17600
rect 13678 17599 13703 17600
rect 13714 17599 13781 17600
rect 13792 17599 13817 17600
rect 13856 17528 13857 17543
rect 13591 17482 13600 17499
rect 13591 17481 13617 17482
rect 12317 17376 12318 17391
rect 12740 17383 12745 17399
rect 12723 17366 12728 17382
rect 13011 17376 13012 17391
rect 13871 17376 13872 17391
rect 13833 17355 13834 17363
rect 13402 17346 13468 17347
rect 13558 17346 13624 17347
rect 13714 17346 13780 17347
rect 13419 17329 13451 17330
rect 13575 17329 13607 17330
rect 13731 17329 13763 17330
rect 12213 17304 12230 17321
rect 12331 17304 12348 17321
rect 12907 17304 12924 17321
rect 13025 17304 13042 17321
rect 13280 17304 13297 17321
rect 13349 17304 13366 17321
rect 13427 17304 13444 17321
rect 13505 17304 13522 17321
rect 13583 17304 13600 17321
rect 13661 17304 13678 17321
rect 13739 17304 13756 17321
rect 13817 17304 13834 17321
rect 13885 17304 13902 17321
rect 12586 17284 12603 17301
rect 12645 17284 12662 17301
rect 14531 17248 14569 17259
rect 31691 17248 31729 17259
rect 12078 17247 12205 17248
rect 12238 17247 12381 17248
rect 12414 17247 12578 17248
rect 12611 17247 12695 17248
rect 12728 17247 12764 17248
rect 12781 17247 12899 17248
rect 12932 17247 13075 17248
rect 13108 17247 13272 17248
rect 13305 17247 13419 17248
rect 13451 17247 13575 17248
rect 13607 17247 13731 17248
rect 13763 17247 13877 17248
rect 13910 17247 13935 17248
rect 13968 17247 13997 17248
rect 12796 17225 12797 17247
rect 12839 17225 12840 17247
rect 14441 17230 14458 17248
rect 14534 17230 14551 17248
rect 14605 17230 14622 17248
rect 14701 17230 14718 17248
rect 14794 17230 14811 17248
rect 14865 17230 14882 17248
rect 14961 17230 14978 17248
rect 15054 17230 15071 17248
rect 15125 17230 15142 17248
rect 15221 17230 15238 17248
rect 31081 17230 31098 17248
rect 31174 17230 31191 17248
rect 31245 17230 31262 17248
rect 31341 17230 31358 17248
rect 31434 17230 31451 17248
rect 31505 17230 31522 17248
rect 31601 17230 31618 17248
rect 31694 17230 31711 17248
rect 31765 17230 31782 17248
rect 12796 17224 12840 17225
rect 14531 17219 14569 17230
rect 31691 17219 31729 17230
rect 12586 17177 12603 17194
rect 12645 17186 12662 17194
rect 12632 17185 12676 17186
rect 12213 17157 12230 17174
rect 12331 17157 12348 17174
rect 12632 17163 12633 17185
rect 12645 17177 12662 17185
rect 12675 17163 12676 17185
rect 31738 17185 31782 17186
rect 12907 17157 12924 17174
rect 13025 17157 13042 17174
rect 13280 17157 13297 17174
rect 13349 17157 13366 17174
rect 13427 17157 13444 17174
rect 13505 17157 13522 17174
rect 13583 17157 13600 17174
rect 13661 17157 13678 17174
rect 13739 17157 13756 17174
rect 13817 17157 13834 17174
rect 13885 17157 13902 17174
rect 31738 17163 31739 17185
rect 31781 17163 31782 17185
rect 13419 17148 13451 17149
rect 13575 17148 13607 17149
rect 13731 17148 13763 17149
rect 13816 17132 13817 17140
rect 13402 17131 13468 17132
rect 13558 17131 13624 17132
rect 13714 17131 13780 17132
rect 12302 17102 12303 17117
rect 12723 17096 12728 17113
rect 12996 17102 12997 17117
rect 13856 17102 13857 17117
rect 12740 17079 12745 17096
rect 13591 17014 13600 17031
rect 13591 17013 13617 17014
rect 13871 16950 13872 16965
rect 13833 16887 13834 16895
rect 12317 16866 12318 16881
rect 13011 16866 13012 16881
rect 13366 16878 13391 16879
rect 13402 16878 13469 16879
rect 13480 16878 13505 16879
rect 13522 16878 13547 16879
rect 13558 16878 13625 16879
rect 13636 16878 13661 16879
rect 13678 16878 13703 16879
rect 13714 16878 13781 16879
rect 13792 16878 13817 16879
rect 12357 16861 12365 16862
rect 13051 16861 13059 16862
rect 13366 16861 13374 16862
rect 13419 16861 13452 16862
rect 13497 16861 13505 16862
rect 13522 16861 13530 16862
rect 13575 16861 13608 16862
rect 13653 16861 13661 16862
rect 13678 16861 13686 16862
rect 13731 16861 13764 16862
rect 13809 16861 13817 16862
rect 12364 16844 12374 16845
rect 12381 16827 12391 16845
rect 13058 16844 13068 16845
rect 13075 16827 13085 16845
rect 13280 16837 13297 16854
rect 13349 16837 13366 16854
rect 13427 16837 13444 16854
rect 13505 16837 13522 16854
rect 13583 16837 13600 16854
rect 13661 16837 13678 16854
rect 13739 16837 13756 16854
rect 13817 16837 13834 16854
rect 13885 16837 13902 16854
rect 12213 16795 12230 16812
rect 12272 16795 12289 16812
rect 12331 16795 12348 16812
rect 12586 16795 12603 16812
rect 12645 16795 12662 16812
rect 12907 16795 12924 16812
rect 12966 16795 12983 16812
rect 13025 16795 13042 16812
rect 12244 16740 12259 16741
rect 12303 16740 12318 16741
rect 12617 16740 12632 16741
rect 12938 16740 12953 16741
rect 12997 16740 13012 16741
rect 13311 16740 13326 16741
rect 13389 16740 13404 16741
rect 13467 16740 13482 16741
rect 13545 16740 13560 16741
rect 13623 16740 13638 16741
rect 13701 16740 13716 16741
rect 13779 16740 13794 16741
rect 13857 16740 13872 16741
rect 12755 16738 12765 16739
rect 12772 16738 12782 16739
rect 14456 16721 14473 16739
rect 14531 16709 14569 16751
rect 14581 16721 14598 16739
rect 14631 16721 14648 16739
rect 14716 16721 14733 16739
rect 14794 16721 14811 16739
rect 14841 16721 14858 16739
rect 14891 16721 14908 16739
rect 14976 16721 14993 16739
rect 15054 16721 15071 16739
rect 15101 16721 15118 16739
rect 15151 16721 15168 16739
rect 15236 16721 15253 16739
rect 31022 16721 31028 16739
rect 31096 16721 31113 16739
rect 31174 16721 31191 16739
rect 31221 16721 31238 16739
rect 31271 16721 31288 16739
rect 31356 16721 31373 16739
rect 31434 16721 31451 16739
rect 31481 16721 31498 16739
rect 31531 16721 31548 16739
rect 31616 16721 31633 16739
rect 31691 16709 31729 16751
rect 31741 16721 31758 16739
rect 31791 16721 31808 16739
rect 12213 16648 12230 16665
rect 12272 16648 12289 16665
rect 12331 16648 12348 16665
rect 12586 16648 12603 16665
rect 12645 16648 12662 16665
rect 12907 16648 12924 16665
rect 12966 16648 12983 16665
rect 13025 16648 13042 16665
rect 12381 16616 12391 16633
rect 13075 16616 13085 16633
rect 12364 16615 12391 16616
rect 13058 16615 13085 16616
rect 12302 16594 12303 16609
rect 12996 16594 12997 16609
rect 13280 16606 13297 16623
rect 13349 16606 13366 16623
rect 13427 16606 13444 16623
rect 13505 16606 13522 16623
rect 13583 16606 13600 16623
rect 13661 16606 13678 16623
rect 13739 16606 13756 16623
rect 13817 16606 13834 16623
rect 13885 16606 13902 16623
rect 13366 16598 13374 16599
rect 13419 16598 13452 16599
rect 13497 16598 13505 16599
rect 13522 16598 13530 16599
rect 13575 16598 13608 16599
rect 13653 16598 13661 16599
rect 13678 16598 13686 16599
rect 13731 16598 13764 16599
rect 13809 16598 13817 16599
rect 13816 16582 13817 16590
rect 13366 16581 13391 16582
rect 13402 16581 13469 16582
rect 13480 16581 13505 16582
rect 13522 16581 13547 16582
rect 13558 16581 13625 16582
rect 13636 16581 13661 16582
rect 13678 16581 13703 16582
rect 13714 16581 13781 16582
rect 13792 16581 13817 16582
rect 13856 16510 13857 16525
rect 13591 16464 13600 16481
rect 13591 16463 13617 16464
rect 12317 16358 12318 16373
rect 12740 16365 12745 16381
rect 12723 16348 12728 16364
rect 13011 16358 13012 16373
rect 13871 16358 13872 16373
rect 13833 16337 13834 16345
rect 13402 16328 13468 16329
rect 13558 16328 13624 16329
rect 13714 16328 13780 16329
rect 13419 16311 13451 16312
rect 13575 16311 13607 16312
rect 13731 16311 13763 16312
rect 12213 16286 12230 16303
rect 12331 16286 12348 16303
rect 12907 16286 12924 16303
rect 13025 16286 13042 16303
rect 13280 16286 13297 16303
rect 13349 16286 13366 16303
rect 13427 16286 13444 16303
rect 13505 16286 13522 16303
rect 13583 16286 13600 16303
rect 13661 16286 13678 16303
rect 13739 16286 13756 16303
rect 13817 16286 13834 16303
rect 13885 16286 13902 16303
rect 12586 16266 12603 16283
rect 12645 16266 12662 16283
rect 14026 16241 14027 16263
rect 14069 16241 14070 16263
rect 14026 16240 14070 16241
rect 14531 16230 14569 16241
rect 31691 16230 31729 16241
rect 12078 16229 12205 16230
rect 12238 16229 12381 16230
rect 12414 16229 12578 16230
rect 12611 16229 12695 16230
rect 12728 16229 12764 16230
rect 12781 16229 12899 16230
rect 12932 16229 13075 16230
rect 13108 16229 13272 16230
rect 13305 16229 13419 16230
rect 13451 16229 13575 16230
rect 13607 16229 13731 16230
rect 13763 16229 13877 16230
rect 13910 16229 13935 16230
rect 13968 16229 13997 16230
rect 14441 16212 14458 16230
rect 14534 16212 14551 16230
rect 14605 16212 14622 16230
rect 14701 16212 14718 16230
rect 14794 16212 14811 16230
rect 14865 16212 14882 16230
rect 14961 16212 14978 16230
rect 15054 16212 15071 16230
rect 15125 16212 15142 16230
rect 15221 16212 15238 16230
rect 31081 16212 31098 16230
rect 31174 16212 31191 16230
rect 31245 16212 31262 16230
rect 31341 16212 31358 16230
rect 31434 16212 31451 16230
rect 31505 16212 31522 16230
rect 31601 16212 31618 16230
rect 31694 16212 31711 16230
rect 31765 16212 31782 16230
rect 8122 16201 8166 16202
rect 8122 16179 8123 16201
rect 8165 16179 8166 16201
rect 12878 16201 12922 16202
rect 14531 16201 14569 16212
rect 31691 16201 31729 16212
rect 31738 16201 31782 16202
rect 12878 16179 12879 16201
rect 12921 16179 12922 16201
rect 31738 16179 31739 16201
rect 31781 16179 31782 16201
rect 12586 16159 12603 16176
rect 12645 16159 12662 16176
rect 12213 16139 12230 16156
rect 12331 16139 12348 16156
rect 12907 16139 12924 16156
rect 13025 16139 13042 16156
rect 13280 16139 13297 16156
rect 13349 16139 13366 16156
rect 13427 16139 13444 16156
rect 13505 16139 13522 16156
rect 13583 16139 13600 16156
rect 13661 16139 13678 16156
rect 13739 16139 13756 16156
rect 13817 16139 13834 16156
rect 13885 16139 13902 16156
rect 13419 16130 13451 16131
rect 13575 16130 13607 16131
rect 13731 16130 13763 16131
rect 13816 16114 13817 16122
rect 13402 16113 13468 16114
rect 13558 16113 13624 16114
rect 13714 16113 13780 16114
rect 12302 16084 12303 16099
rect 12723 16078 12728 16095
rect 12996 16084 12997 16099
rect 13856 16084 13857 16099
rect 12740 16061 12745 16078
rect 13591 15996 13600 16013
rect 13591 15995 13617 15996
rect 13871 15932 13872 15947
rect 13833 15869 13834 15877
rect 12317 15848 12318 15863
rect 13011 15848 13012 15863
rect 13366 15860 13391 15861
rect 13402 15860 13469 15861
rect 13480 15860 13505 15861
rect 13522 15860 13547 15861
rect 13558 15860 13625 15861
rect 13636 15860 13661 15861
rect 13678 15860 13703 15861
rect 13714 15860 13781 15861
rect 13792 15860 13817 15861
rect 12357 15843 12365 15844
rect 13051 15843 13059 15844
rect 13366 15843 13374 15844
rect 13419 15843 13452 15844
rect 13497 15843 13505 15844
rect 13522 15843 13530 15844
rect 13575 15843 13608 15844
rect 13653 15843 13661 15844
rect 13678 15843 13686 15844
rect 13731 15843 13764 15844
rect 13809 15843 13817 15844
rect 7494 15798 7511 15820
rect 7554 15798 7571 15820
rect 7637 15798 7654 15820
rect 7697 15798 7714 15820
rect 7741 15798 7758 15820
rect 7801 15798 7818 15820
rect 7852 15798 7869 15820
rect 7988 15798 8005 15820
rect 8037 15798 8054 15820
rect 8095 15787 8133 15831
rect 12364 15826 12374 15827
rect 8217 15798 8234 15820
rect 8277 15798 8294 15820
rect 8321 15798 8338 15820
rect 8381 15798 8398 15820
rect 8432 15798 8449 15820
rect 8592 15798 8609 15820
rect 8641 15798 8658 15820
rect 8701 15798 8718 15820
rect 12381 15809 12391 15827
rect 13058 15826 13068 15827
rect 13075 15809 13085 15827
rect 13280 15819 13297 15836
rect 13349 15819 13366 15836
rect 13427 15819 13444 15836
rect 13505 15819 13522 15836
rect 13583 15819 13600 15836
rect 13661 15819 13678 15836
rect 13739 15819 13756 15836
rect 13817 15819 13834 15836
rect 13885 15819 13902 15836
rect 12213 15777 12230 15794
rect 12272 15777 12289 15794
rect 12331 15777 12348 15794
rect 12586 15777 12603 15794
rect 12645 15777 12662 15794
rect 12907 15777 12924 15794
rect 12966 15777 12983 15794
rect 13025 15777 13042 15794
rect 12796 15749 12797 15771
rect 12839 15749 12840 15771
rect 12796 15748 12840 15749
rect 13944 15749 13945 15771
rect 13987 15749 13988 15771
rect 13944 15748 13988 15749
rect 12244 15722 12259 15723
rect 12303 15722 12318 15723
rect 12617 15722 12632 15723
rect 12938 15722 12953 15723
rect 12997 15722 13012 15723
rect 13311 15722 13326 15723
rect 13389 15722 13404 15723
rect 13467 15722 13482 15723
rect 13545 15722 13560 15723
rect 13623 15722 13638 15723
rect 13701 15722 13716 15723
rect 13779 15722 13794 15723
rect 13857 15722 13872 15723
rect 12755 15720 12765 15721
rect 12772 15720 12782 15721
rect 12714 15709 12758 15710
rect 12714 15687 12715 15709
rect 12757 15687 12758 15709
rect 14456 15703 14473 15721
rect 14531 15691 14569 15733
rect 14581 15703 14598 15721
rect 14631 15710 14648 15721
rect 14600 15709 14648 15710
rect 14600 15687 14601 15709
rect 14631 15703 14648 15709
rect 14716 15703 14733 15721
rect 14794 15703 14811 15721
rect 14841 15703 14858 15721
rect 14891 15703 14908 15721
rect 14976 15703 14993 15721
rect 15054 15703 15071 15721
rect 15101 15703 15118 15721
rect 15151 15703 15168 15721
rect 15236 15703 15253 15721
rect 31022 15703 31028 15721
rect 31096 15703 31113 15721
rect 31174 15703 31191 15721
rect 31221 15703 31238 15721
rect 31271 15703 31288 15721
rect 31356 15703 31373 15721
rect 31434 15703 31451 15721
rect 31481 15703 31498 15721
rect 31531 15703 31548 15721
rect 31616 15703 31633 15721
rect 14643 15687 14644 15703
rect 31691 15691 31729 15733
rect 31741 15703 31758 15721
rect 31791 15703 31808 15721
rect 12213 15630 12230 15647
rect 12272 15630 12289 15647
rect 12331 15630 12348 15647
rect 12586 15630 12603 15647
rect 12645 15630 12662 15647
rect 12907 15630 12924 15647
rect 12966 15630 12983 15647
rect 13025 15630 13042 15647
rect 12381 15598 12391 15615
rect 13075 15598 13085 15615
rect 12364 15597 12391 15598
rect 13058 15597 13085 15598
rect 12302 15576 12303 15591
rect 12996 15576 12997 15591
rect 13280 15588 13297 15605
rect 13349 15588 13366 15605
rect 13427 15588 13444 15605
rect 13505 15588 13522 15605
rect 13583 15588 13600 15605
rect 13661 15588 13678 15605
rect 13739 15588 13756 15605
rect 13817 15588 13834 15605
rect 13885 15588 13902 15605
rect 13366 15580 13374 15581
rect 13419 15580 13452 15581
rect 13497 15580 13505 15581
rect 13522 15580 13530 15581
rect 13575 15580 13608 15581
rect 13653 15580 13661 15581
rect 13678 15580 13686 15581
rect 13731 15580 13764 15581
rect 13809 15580 13817 15581
rect 13816 15564 13817 15572
rect 13366 15563 13391 15564
rect 13402 15563 13469 15564
rect 13480 15563 13505 15564
rect 13522 15563 13547 15564
rect 13558 15563 13625 15564
rect 13636 15563 13661 15564
rect 13678 15563 13703 15564
rect 13714 15563 13781 15564
rect 13792 15563 13817 15564
rect 13856 15492 13857 15507
rect 13591 15446 13600 15463
rect 13591 15445 13617 15446
rect 8095 15412 8133 15423
rect 7515 15394 7532 15412
rect 7589 15394 7606 15412
rect 7658 15394 7675 15412
rect 7737 15394 7754 15412
rect 7810 15394 7827 15412
rect 7965 15394 7982 15412
rect 8044 15394 8061 15412
rect 8123 15394 8140 15412
rect 8238 15394 8255 15412
rect 8317 15394 8334 15412
rect 8390 15394 8407 15412
rect 8569 15394 8586 15412
rect 8648 15394 8665 15412
rect 8095 15383 8133 15394
rect 8040 15381 8084 15382
rect 8040 15359 8041 15381
rect 8083 15359 8084 15381
rect 12317 15340 12318 15355
rect 12740 15347 12745 15363
rect 12723 15330 12728 15346
rect 13011 15340 13012 15355
rect 13871 15340 13872 15355
rect 13833 15319 13834 15327
rect 13402 15310 13468 15311
rect 13558 15310 13624 15311
rect 13714 15310 13780 15311
rect 13419 15293 13451 15294
rect 13575 15293 13607 15294
rect 13731 15293 13763 15294
rect 12213 15268 12230 15285
rect 12331 15268 12348 15285
rect 12907 15268 12924 15285
rect 13025 15268 13042 15285
rect 13280 15268 13297 15285
rect 13349 15268 13366 15285
rect 13427 15268 13444 15285
rect 13505 15268 13522 15285
rect 13583 15268 13600 15285
rect 13661 15268 13678 15285
rect 13739 15268 13756 15285
rect 13817 15268 13834 15285
rect 13885 15268 13902 15285
rect 12586 15248 12603 15265
rect 12645 15248 12662 15265
rect 14026 15257 14027 15279
rect 14069 15257 14070 15279
rect 14026 15256 14070 15257
rect 14531 15212 14569 15223
rect 31691 15212 31729 15223
rect 12078 15211 12205 15212
rect 12238 15211 12381 15212
rect 12414 15211 12578 15212
rect 12611 15211 12695 15212
rect 12728 15211 12764 15212
rect 12781 15211 12899 15212
rect 12932 15211 13075 15212
rect 13108 15211 13272 15212
rect 13305 15211 13419 15212
rect 13451 15211 13575 15212
rect 13607 15211 13731 15212
rect 13763 15211 13877 15212
rect 13910 15211 13935 15212
rect 13968 15211 13997 15212
rect 14441 15194 14458 15212
rect 14534 15194 14551 15212
rect 14605 15194 14622 15212
rect 14701 15194 14718 15212
rect 14794 15194 14811 15212
rect 14865 15194 14882 15212
rect 14961 15194 14978 15212
rect 15054 15194 15071 15212
rect 15125 15194 15142 15212
rect 15221 15194 15238 15212
rect 31081 15194 31098 15212
rect 31174 15194 31191 15212
rect 31245 15194 31262 15212
rect 31341 15194 31358 15212
rect 31434 15194 31451 15212
rect 31505 15194 31522 15212
rect 31601 15194 31618 15212
rect 31694 15194 31711 15212
rect 31765 15194 31782 15212
rect 14531 15183 14569 15194
rect 31691 15183 31729 15194
rect 12586 15141 12603 15158
rect 12645 15141 12662 15158
rect 12213 15121 12230 15138
rect 12331 15121 12348 15138
rect 12907 15121 12924 15138
rect 13025 15121 13042 15138
rect 13280 15121 13297 15138
rect 13349 15121 13366 15138
rect 13427 15121 13444 15138
rect 13505 15121 13522 15138
rect 13583 15121 13600 15138
rect 13661 15121 13678 15138
rect 13739 15121 13756 15138
rect 13817 15121 13834 15138
rect 13885 15121 13902 15138
rect 13419 15112 13451 15113
rect 13575 15112 13607 15113
rect 13731 15112 13763 15113
rect 13816 15096 13817 15104
rect 13402 15095 13468 15096
rect 13558 15095 13624 15096
rect 13714 15095 13780 15096
rect 12302 15066 12303 15081
rect 12723 15060 12728 15077
rect 12996 15066 12997 15081
rect 13856 15066 13857 15081
rect 12740 15043 12745 15060
rect 7958 15011 7959 15033
rect 8001 15011 8002 15033
rect 7958 15010 8002 15011
rect 7494 14986 7511 15008
rect 7554 14986 7571 15008
rect 7637 14986 7654 15008
rect 7697 14986 7714 15008
rect 7741 14986 7758 15008
rect 7801 14986 7818 15008
rect 7852 14986 7869 15008
rect 7988 14986 8005 15008
rect 8037 14986 8054 15008
rect 8095 14975 8133 15019
rect 8217 14986 8234 15008
rect 8277 14986 8294 15008
rect 8321 14986 8338 15008
rect 8381 14986 8398 15008
rect 8432 14986 8449 15008
rect 8592 14986 8609 15008
rect 8641 14986 8658 15008
rect 8701 14986 8718 15008
rect 13591 14978 13600 14995
rect 13591 14977 13617 14978
rect 8122 14971 8166 14972
rect 8122 14949 8123 14971
rect 8165 14949 8166 14971
rect 13871 14914 13872 14929
rect 13833 14851 13834 14859
rect 12317 14830 12318 14845
rect 13011 14830 13012 14845
rect 13366 14842 13391 14843
rect 13402 14842 13469 14843
rect 13480 14842 13505 14843
rect 13522 14842 13547 14843
rect 13558 14842 13625 14843
rect 13636 14842 13661 14843
rect 13678 14842 13703 14843
rect 13714 14842 13781 14843
rect 13792 14842 13817 14843
rect 12357 14825 12365 14826
rect 13051 14825 13059 14826
rect 13366 14825 13374 14826
rect 13419 14825 13452 14826
rect 13497 14825 13505 14826
rect 13522 14825 13530 14826
rect 13575 14825 13608 14826
rect 13653 14825 13661 14826
rect 13678 14825 13686 14826
rect 13731 14825 13764 14826
rect 13809 14825 13817 14826
rect 12364 14808 12374 14809
rect 12381 14791 12391 14809
rect 13058 14808 13068 14809
rect 13075 14791 13085 14809
rect 13280 14801 13297 14818
rect 13349 14801 13366 14818
rect 13427 14801 13444 14818
rect 13505 14801 13522 14818
rect 13583 14801 13600 14818
rect 13661 14801 13678 14818
rect 13739 14801 13756 14818
rect 13817 14801 13834 14818
rect 13885 14801 13902 14818
rect 12213 14759 12230 14776
rect 12272 14759 12289 14776
rect 12331 14759 12348 14776
rect 12586 14759 12603 14776
rect 12645 14759 12662 14776
rect 12907 14759 12924 14776
rect 12966 14759 12983 14776
rect 13025 14759 13042 14776
rect 12244 14704 12259 14705
rect 12303 14704 12318 14705
rect 12617 14704 12632 14705
rect 12938 14704 12953 14705
rect 12997 14704 13012 14705
rect 13311 14704 13326 14705
rect 13389 14704 13404 14705
rect 13467 14704 13482 14705
rect 13545 14704 13560 14705
rect 13623 14704 13638 14705
rect 13701 14704 13716 14705
rect 13779 14704 13794 14705
rect 13857 14704 13872 14705
rect 12755 14702 12765 14703
rect 12772 14702 12782 14703
rect 14456 14685 14473 14703
rect 14531 14673 14569 14715
rect 14581 14685 14598 14703
rect 14631 14685 14648 14703
rect 14716 14685 14733 14703
rect 14794 14685 14811 14703
rect 14841 14685 14858 14703
rect 14891 14685 14908 14703
rect 14976 14685 14993 14703
rect 15054 14685 15071 14703
rect 15101 14685 15118 14703
rect 15151 14685 15168 14703
rect 15236 14685 15253 14703
rect 31022 14685 31028 14703
rect 31096 14685 31113 14703
rect 31174 14685 31191 14703
rect 31221 14685 31238 14703
rect 31271 14685 31288 14703
rect 31356 14685 31373 14703
rect 31434 14685 31451 14703
rect 31481 14685 31498 14703
rect 31531 14685 31548 14703
rect 31616 14685 31633 14703
rect 31691 14673 31729 14715
rect 31741 14685 31758 14703
rect 31791 14685 31808 14703
rect 12714 14643 12758 14644
rect 12213 14612 12230 14629
rect 12272 14612 12289 14629
rect 12331 14612 12348 14629
rect 12586 14612 12603 14629
rect 12645 14612 12662 14629
rect 12714 14621 12715 14643
rect 12757 14621 12758 14643
rect 12907 14612 12924 14629
rect 12966 14612 12983 14629
rect 13025 14612 13042 14629
rect 8095 14600 8133 14611
rect 7515 14582 7532 14600
rect 7589 14582 7606 14600
rect 7658 14582 7675 14600
rect 7737 14582 7754 14600
rect 7810 14582 7827 14600
rect 7965 14582 7982 14600
rect 8044 14582 8061 14600
rect 8123 14582 8140 14600
rect 8238 14582 8255 14600
rect 8317 14582 8334 14600
rect 8390 14582 8407 14600
rect 8569 14582 8586 14600
rect 8648 14582 8665 14600
rect 8095 14571 8133 14582
rect 12381 14580 12391 14597
rect 13075 14580 13085 14597
rect 12364 14579 12391 14580
rect 13058 14579 13085 14580
rect 9516 14561 9560 14562
rect 9516 14539 9517 14561
rect 9559 14539 9560 14561
rect 12302 14558 12303 14573
rect 12996 14558 12997 14573
rect 13280 14570 13297 14587
rect 13349 14570 13366 14587
rect 13427 14570 13444 14587
rect 13505 14570 13522 14587
rect 13583 14570 13600 14587
rect 13661 14570 13678 14587
rect 13739 14570 13756 14587
rect 13817 14570 13834 14587
rect 13885 14570 13902 14587
rect 13366 14562 13374 14563
rect 13419 14562 13452 14563
rect 13497 14562 13505 14563
rect 13522 14562 13530 14563
rect 13575 14562 13608 14563
rect 13653 14562 13661 14563
rect 13678 14562 13686 14563
rect 13731 14562 13764 14563
rect 13809 14562 13817 14563
rect 13816 14546 13817 14554
rect 13366 14545 13391 14546
rect 13402 14545 13469 14546
rect 13480 14545 13505 14546
rect 13522 14545 13547 14546
rect 13558 14545 13625 14546
rect 13636 14545 13661 14546
rect 13678 14545 13703 14546
rect 13714 14545 13781 14546
rect 13792 14545 13817 14546
rect 13856 14474 13857 14489
rect 13591 14428 13600 14445
rect 13591 14427 13617 14428
rect 7593 14406 7645 14424
rect 7517 14397 7561 14401
rect 7517 14361 7521 14397
rect 7555 14361 7561 14397
rect 7585 14376 7675 14394
rect 7585 14364 7591 14376
rect 7517 14357 7561 14361
rect 12317 14322 12318 14337
rect 12740 14329 12745 14345
rect 12723 14312 12728 14328
rect 13011 14322 13012 14337
rect 13871 14322 13872 14337
rect 13833 14301 13834 14309
rect 13402 14292 13468 14293
rect 13558 14292 13624 14293
rect 13714 14292 13780 14293
rect 13419 14275 13451 14276
rect 13575 14275 13607 14276
rect 13731 14275 13763 14276
rect 12213 14250 12230 14267
rect 12331 14250 12348 14267
rect 12907 14250 12924 14267
rect 13025 14250 13042 14267
rect 13280 14250 13297 14267
rect 13349 14250 13366 14267
rect 13427 14250 13444 14267
rect 13505 14250 13522 14267
rect 13583 14250 13600 14267
rect 13661 14250 13678 14267
rect 13739 14250 13756 14267
rect 13817 14250 13834 14267
rect 13885 14250 13902 14267
rect 12586 14230 12603 14247
rect 12645 14230 12662 14247
rect 12796 14194 12797 14213
rect 12839 14194 12840 14213
rect 12078 14193 12205 14194
rect 12238 14193 12381 14194
rect 12414 14193 12578 14194
rect 12611 14193 12695 14194
rect 12728 14193 12764 14194
rect 12781 14193 12899 14194
rect 12932 14193 13075 14194
rect 13108 14193 13272 14194
rect 13305 14193 13419 14194
rect 13451 14193 13575 14194
rect 13607 14193 13731 14194
rect 13763 14193 13877 14194
rect 13910 14193 13935 14194
rect 13968 14193 13997 14194
rect 12796 14191 12797 14193
rect 12839 14191 12840 14193
rect 12796 14190 12840 14191
rect 14026 14191 14027 14213
rect 14069 14191 14070 14213
rect 14531 14194 14569 14205
rect 31691 14194 31729 14205
rect 14026 14190 14070 14191
rect 14441 14176 14458 14194
rect 14534 14176 14551 14194
rect 14605 14176 14622 14194
rect 14701 14176 14718 14194
rect 14794 14176 14811 14194
rect 14865 14176 14882 14194
rect 14961 14176 14978 14194
rect 15054 14176 15071 14194
rect 15125 14176 15142 14194
rect 15221 14176 15238 14194
rect 31081 14176 31098 14194
rect 31174 14176 31191 14194
rect 31245 14176 31262 14194
rect 31341 14176 31358 14194
rect 31434 14176 31451 14194
rect 31505 14176 31522 14194
rect 31601 14176 31618 14194
rect 31694 14176 31711 14194
rect 31765 14176 31782 14194
rect 14531 14165 14569 14176
rect 31691 14165 31729 14176
rect 12796 14151 12840 14152
rect 11041 14123 11058 14140
rect 11100 14123 11117 14140
rect 12586 14123 12603 14140
rect 12645 14123 12662 14140
rect 12796 14129 12797 14151
rect 12839 14129 12840 14151
rect 14600 14151 14644 14152
rect 14600 14129 14601 14151
rect 14643 14129 14644 14151
rect 31656 14151 31700 14152
rect 31656 14129 31657 14151
rect 31699 14129 31700 14151
rect 10549 14103 10566 14120
rect 10726 14103 10743 14120
rect 12213 14103 12230 14120
rect 12331 14103 12348 14120
rect 12907 14103 12924 14120
rect 13025 14103 13042 14120
rect 13280 14103 13297 14120
rect 13349 14103 13366 14120
rect 13427 14103 13444 14120
rect 13505 14103 13522 14120
rect 13583 14103 13600 14120
rect 13661 14103 13678 14120
rect 13739 14103 13756 14120
rect 13817 14103 13834 14120
rect 13885 14103 13902 14120
rect 13419 14094 13451 14095
rect 13575 14094 13607 14095
rect 13731 14094 13763 14095
rect 13816 14078 13817 14086
rect 13402 14077 13468 14078
rect 13558 14077 13624 14078
rect 13714 14077 13780 14078
rect 10638 14048 10639 14063
rect 12302 14048 12303 14063
rect 12723 14042 12728 14059
rect 12996 14048 12997 14063
rect 13856 14048 13857 14063
rect 12740 14025 12745 14042
rect 11101 13950 11117 13967
rect 13591 13960 13600 13977
rect 13591 13959 13617 13960
rect 11101 13949 11134 13950
rect 10743 13852 10751 13885
rect 10760 13835 10768 13902
rect 13871 13896 13872 13911
rect 13833 13833 13834 13841
rect 10653 13812 10654 13827
rect 12317 13812 12318 13827
rect 13011 13812 13012 13827
rect 13366 13824 13391 13825
rect 13402 13824 13469 13825
rect 13480 13824 13505 13825
rect 13522 13824 13547 13825
rect 13558 13824 13625 13825
rect 13636 13824 13661 13825
rect 13678 13824 13703 13825
rect 13714 13824 13781 13825
rect 13792 13824 13817 13825
rect 12357 13807 12365 13808
rect 13051 13807 13059 13808
rect 13366 13807 13374 13808
rect 13419 13807 13452 13808
rect 13497 13807 13505 13808
rect 13522 13807 13530 13808
rect 13575 13807 13608 13808
rect 13653 13807 13661 13808
rect 13678 13807 13686 13808
rect 13731 13807 13764 13808
rect 13809 13807 13817 13808
rect 10751 13799 10760 13800
rect 12364 13790 12374 13791
rect 10625 13782 10726 13783
rect 10743 13782 10768 13783
rect 12381 13773 12391 13791
rect 13058 13790 13068 13791
rect 13075 13773 13085 13791
rect 13280 13783 13297 13800
rect 13349 13783 13366 13800
rect 13427 13783 13444 13800
rect 13505 13783 13522 13800
rect 13583 13783 13600 13800
rect 13661 13783 13678 13800
rect 13739 13783 13756 13800
rect 13817 13783 13834 13800
rect 13885 13783 13902 13800
rect 10625 13765 10633 13766
rect 10659 13765 10692 13766
rect 10718 13765 10726 13766
rect 10743 13765 10751 13766
rect 10549 13741 10566 13758
rect 10608 13741 10625 13758
rect 10667 13741 10684 13758
rect 10726 13741 10743 13758
rect 11041 13741 11058 13758
rect 11100 13741 11117 13758
rect 12213 13741 12230 13758
rect 12272 13741 12289 13758
rect 12331 13741 12348 13758
rect 12586 13741 12603 13758
rect 12645 13741 12662 13758
rect 12907 13741 12924 13758
rect 12966 13741 12983 13758
rect 13025 13741 13042 13758
rect 13944 13699 13945 13721
rect 13987 13699 13988 13721
rect 13944 13698 13988 13699
rect 10580 13686 10595 13687
rect 10639 13686 10654 13687
rect 10698 13686 10713 13687
rect 11072 13686 11087 13687
rect 12244 13686 12259 13687
rect 12303 13686 12318 13687
rect 12617 13686 12632 13687
rect 12938 13686 12953 13687
rect 12997 13686 13012 13687
rect 13311 13686 13326 13687
rect 13389 13686 13404 13687
rect 13467 13686 13482 13687
rect 13545 13686 13560 13687
rect 13623 13686 13638 13687
rect 13701 13686 13716 13687
rect 13779 13686 13794 13687
rect 13857 13686 13872 13687
rect 12755 13684 12765 13685
rect 12772 13684 12782 13685
rect 14456 13667 14473 13685
rect 14531 13655 14569 13697
rect 14581 13667 14598 13685
rect 14631 13667 14648 13685
rect 14716 13667 14733 13685
rect 14794 13667 14811 13685
rect 14841 13667 14858 13685
rect 14891 13667 14908 13685
rect 14976 13667 14993 13685
rect 15054 13667 15071 13685
rect 15101 13667 15118 13685
rect 15151 13667 15168 13685
rect 15236 13667 15253 13685
rect 31022 13667 31028 13685
rect 31096 13667 31113 13685
rect 31174 13667 31191 13685
rect 31221 13667 31238 13685
rect 31271 13667 31288 13685
rect 31356 13667 31373 13685
rect 31434 13667 31451 13685
rect 31481 13667 31498 13685
rect 31531 13667 31548 13685
rect 31616 13667 31633 13685
rect 31691 13655 31729 13697
rect 31741 13667 31758 13685
rect 31791 13667 31808 13685
rect 10549 13594 10566 13611
rect 10608 13594 10625 13611
rect 10667 13594 10684 13611
rect 10726 13594 10743 13611
rect 11041 13594 11058 13611
rect 11100 13594 11117 13611
rect 12213 13594 12230 13611
rect 12272 13594 12289 13611
rect 12331 13594 12348 13611
rect 12586 13594 12603 13611
rect 12645 13594 12662 13611
rect 12907 13594 12924 13611
rect 12966 13594 12983 13611
rect 13025 13594 13042 13611
rect 10625 13586 10633 13587
rect 10659 13586 10692 13587
rect 10718 13586 10726 13587
rect 10743 13586 10751 13587
rect 10625 13569 10726 13570
rect 10743 13569 10777 13570
rect 12381 13562 12391 13579
rect 13075 13562 13085 13579
rect 12364 13561 12391 13562
rect 13058 13561 13085 13562
rect 10638 13540 10639 13555
rect 12302 13540 12303 13555
rect 12996 13540 12997 13555
rect 13280 13552 13297 13569
rect 13349 13552 13366 13569
rect 13427 13552 13444 13569
rect 13505 13552 13522 13569
rect 13583 13552 13600 13569
rect 13661 13552 13678 13569
rect 13739 13552 13756 13569
rect 13817 13552 13834 13569
rect 13885 13552 13902 13569
rect 13366 13544 13374 13545
rect 13419 13544 13452 13545
rect 13497 13544 13505 13545
rect 13522 13544 13530 13545
rect 13575 13544 13608 13545
rect 13653 13544 13661 13545
rect 13678 13544 13686 13545
rect 13731 13544 13764 13545
rect 13809 13544 13817 13545
rect 13816 13528 13817 13536
rect 13366 13527 13391 13528
rect 13402 13527 13469 13528
rect 13480 13527 13505 13528
rect 13522 13527 13547 13528
rect 13558 13527 13625 13528
rect 13636 13527 13661 13528
rect 13678 13527 13703 13528
rect 13714 13527 13781 13528
rect 13792 13527 13817 13528
rect 10743 13467 10751 13500
rect 10760 13450 10768 13517
rect 13856 13456 13857 13471
rect 11101 13420 11117 13437
rect 11101 13419 11134 13420
rect 13591 13410 13600 13427
rect 13591 13409 13617 13410
rect 10653 13304 10654 13319
rect 12317 13304 12318 13319
rect 12740 13311 12745 13327
rect 12723 13294 12728 13310
rect 13011 13304 13012 13319
rect 13871 13304 13872 13319
rect 13833 13283 13834 13291
rect 13402 13274 13468 13275
rect 13558 13274 13624 13275
rect 13714 13274 13780 13275
rect 13419 13257 13451 13258
rect 13575 13257 13607 13258
rect 13731 13257 13763 13258
rect 10549 13232 10566 13249
rect 10726 13232 10743 13249
rect 12213 13232 12230 13249
rect 12331 13232 12348 13249
rect 12907 13232 12924 13249
rect 13025 13232 13042 13249
rect 13280 13232 13297 13249
rect 13349 13232 13366 13249
rect 13427 13232 13444 13249
rect 13505 13232 13522 13249
rect 13583 13232 13600 13249
rect 13661 13232 13678 13249
rect 13739 13232 13756 13249
rect 13817 13232 13834 13249
rect 13885 13232 13902 13249
rect 9598 13207 9599 13229
rect 9641 13207 9642 13229
rect 11041 13212 11058 13229
rect 11100 13212 11117 13229
rect 12586 13212 12603 13229
rect 12645 13212 12662 13229
rect 9598 13206 9642 13207
rect 14531 13176 14569 13187
rect 31691 13176 31729 13187
rect 12078 13175 12205 13176
rect 12238 13175 12381 13176
rect 12414 13175 12578 13176
rect 12611 13175 12695 13176
rect 12728 13175 12764 13176
rect 12781 13175 12899 13176
rect 12932 13175 13075 13176
rect 13108 13175 13272 13176
rect 13305 13175 13419 13176
rect 13451 13175 13575 13176
rect 13607 13175 13731 13176
rect 13763 13175 13877 13176
rect 13910 13175 13935 13176
rect 13968 13175 13997 13176
rect 10418 13167 10462 13168
rect 10418 13145 10419 13167
rect 10461 13145 10462 13167
rect 12878 13167 12922 13168
rect 12878 13145 12879 13167
rect 12921 13145 12922 13167
rect 14441 13158 14458 13176
rect 14534 13158 14551 13176
rect 14605 13158 14622 13176
rect 14701 13158 14718 13176
rect 14794 13158 14811 13176
rect 14865 13158 14882 13176
rect 14961 13158 14978 13176
rect 15054 13158 15071 13176
rect 15125 13158 15142 13176
rect 15221 13158 15238 13176
rect 31081 13158 31098 13176
rect 31174 13158 31191 13176
rect 31245 13158 31262 13176
rect 31341 13158 31358 13176
rect 31434 13158 31451 13176
rect 31505 13158 31522 13176
rect 31601 13158 31618 13176
rect 31694 13158 31711 13176
rect 31765 13158 31782 13176
rect 14531 13147 14569 13158
rect 31691 13147 31729 13158
rect 11041 13105 11058 13122
rect 11100 13105 11117 13122
rect 12586 13105 12603 13122
rect 12645 13105 12662 13122
rect 10549 13085 10566 13102
rect 10726 13085 10743 13102
rect 12213 13085 12230 13102
rect 12331 13085 12348 13102
rect 12907 13085 12924 13102
rect 13025 13085 13042 13102
rect 13280 13085 13297 13102
rect 13349 13085 13366 13102
rect 13427 13085 13444 13102
rect 13505 13085 13522 13102
rect 13583 13085 13600 13102
rect 13661 13085 13678 13102
rect 13739 13085 13756 13102
rect 13817 13085 13834 13102
rect 13885 13085 13902 13102
rect 13419 13076 13451 13077
rect 13575 13076 13607 13077
rect 13731 13076 13763 13077
rect 13816 13060 13817 13068
rect 13402 13059 13468 13060
rect 13558 13059 13624 13060
rect 13714 13059 13780 13060
rect 10638 13030 10639 13045
rect 12302 13030 12303 13045
rect 12723 13024 12728 13041
rect 12996 13030 12997 13045
rect 13856 13030 13857 13045
rect 12740 13007 12745 13024
rect 11101 12932 11117 12949
rect 13591 12942 13600 12959
rect 13591 12941 13617 12942
rect 11101 12931 11134 12932
rect 10743 12834 10751 12867
rect 10760 12817 10768 12884
rect 13871 12878 13872 12893
rect 13833 12815 13834 12823
rect 10653 12794 10654 12809
rect 12317 12794 12318 12809
rect 13011 12794 13012 12809
rect 13366 12806 13391 12807
rect 13402 12806 13469 12807
rect 13480 12806 13505 12807
rect 13522 12806 13547 12807
rect 13558 12806 13625 12807
rect 13636 12806 13661 12807
rect 13678 12806 13703 12807
rect 13714 12806 13781 12807
rect 13792 12806 13817 12807
rect 12357 12789 12365 12790
rect 13051 12789 13059 12790
rect 13366 12789 13374 12790
rect 13419 12789 13452 12790
rect 13497 12789 13505 12790
rect 13522 12789 13530 12790
rect 13575 12789 13608 12790
rect 13653 12789 13661 12790
rect 13678 12789 13686 12790
rect 13731 12789 13764 12790
rect 13809 12789 13817 12790
rect 10751 12781 10760 12782
rect 12364 12772 12374 12773
rect 10625 12764 10726 12765
rect 10743 12764 10768 12765
rect 12381 12755 12391 12773
rect 13058 12772 13068 12773
rect 13075 12755 13085 12773
rect 13280 12765 13297 12782
rect 13349 12765 13366 12782
rect 13427 12765 13444 12782
rect 13505 12765 13522 12782
rect 13583 12765 13600 12782
rect 13661 12765 13678 12782
rect 13739 12765 13756 12782
rect 13817 12765 13834 12782
rect 13885 12765 13902 12782
rect 10625 12747 10633 12748
rect 10659 12747 10692 12748
rect 10718 12747 10726 12748
rect 10743 12747 10751 12748
rect 10336 12715 10337 12737
rect 10379 12715 10380 12737
rect 10549 12723 10566 12740
rect 10608 12723 10625 12740
rect 10667 12723 10684 12740
rect 10726 12723 10743 12740
rect 11041 12723 11058 12740
rect 11100 12723 11117 12740
rect 12213 12723 12230 12740
rect 12272 12723 12289 12740
rect 12331 12723 12348 12740
rect 12586 12723 12603 12740
rect 12645 12723 12662 12740
rect 10336 12714 10380 12715
rect 12714 12715 12715 12737
rect 12757 12715 12758 12737
rect 12907 12723 12924 12740
rect 12966 12723 12983 12740
rect 13025 12723 13042 12740
rect 12714 12714 12758 12715
rect 14518 12715 14519 12737
rect 14561 12715 14562 12737
rect 14518 12714 14562 12715
rect 12796 12675 12840 12676
rect 10580 12668 10595 12669
rect 10639 12668 10654 12669
rect 10698 12668 10713 12669
rect 11072 12668 11087 12669
rect 12244 12668 12259 12669
rect 12303 12668 12318 12669
rect 12617 12668 12632 12669
rect 12755 12666 12765 12667
rect 12772 12666 12782 12667
rect 12796 12653 12797 12675
rect 12839 12653 12840 12675
rect 13944 12675 13988 12676
rect 12938 12668 12953 12669
rect 12997 12668 13012 12669
rect 13311 12668 13326 12669
rect 13389 12668 13404 12669
rect 13467 12668 13482 12669
rect 13545 12668 13560 12669
rect 13623 12668 13638 12669
rect 13701 12668 13716 12669
rect 13779 12668 13794 12669
rect 13857 12668 13872 12669
rect 13944 12653 13945 12675
rect 13987 12653 13988 12675
rect 14456 12649 14473 12667
rect 14531 12637 14569 12679
rect 14581 12649 14598 12667
rect 14631 12649 14648 12667
rect 14716 12649 14733 12667
rect 14794 12649 14811 12667
rect 14841 12649 14858 12667
rect 14891 12649 14908 12667
rect 14976 12649 14993 12667
rect 15054 12649 15071 12667
rect 15101 12649 15118 12667
rect 15151 12649 15168 12667
rect 15236 12649 15253 12667
rect 31022 12649 31028 12667
rect 31096 12649 31113 12667
rect 31174 12649 31191 12667
rect 31221 12649 31238 12667
rect 31271 12649 31288 12667
rect 31356 12649 31373 12667
rect 31434 12649 31451 12667
rect 31481 12649 31498 12667
rect 31531 12649 31548 12667
rect 31616 12649 31633 12667
rect 31691 12637 31729 12679
rect 31741 12649 31758 12667
rect 31791 12649 31808 12667
rect 10549 12576 10566 12593
rect 10608 12576 10625 12593
rect 10667 12576 10684 12593
rect 10726 12576 10743 12593
rect 11041 12576 11058 12593
rect 11100 12576 11117 12593
rect 12213 12576 12230 12593
rect 12272 12576 12289 12593
rect 12331 12576 12348 12593
rect 12586 12576 12603 12593
rect 12645 12576 12662 12593
rect 12907 12576 12924 12593
rect 12966 12576 12983 12593
rect 13025 12576 13042 12593
rect 10625 12568 10633 12569
rect 10659 12568 10692 12569
rect 10718 12568 10726 12569
rect 10743 12568 10751 12569
rect 10625 12551 10726 12552
rect 10743 12551 10777 12552
rect 12381 12544 12391 12561
rect 13075 12544 13085 12561
rect 12364 12543 12391 12544
rect 13058 12543 13085 12544
rect 10638 12522 10639 12537
rect 12302 12522 12303 12537
rect 12996 12522 12997 12537
rect 13280 12534 13297 12551
rect 13349 12534 13366 12551
rect 13427 12534 13444 12551
rect 13505 12534 13522 12551
rect 13583 12534 13600 12551
rect 13661 12534 13678 12551
rect 13739 12534 13756 12551
rect 13817 12534 13834 12551
rect 13885 12534 13902 12551
rect 13366 12526 13374 12527
rect 13419 12526 13452 12527
rect 13497 12526 13505 12527
rect 13522 12526 13530 12527
rect 13575 12526 13608 12527
rect 13653 12526 13661 12527
rect 13678 12526 13686 12527
rect 13731 12526 13764 12527
rect 13809 12526 13817 12527
rect 13816 12510 13817 12518
rect 13366 12509 13391 12510
rect 13402 12509 13469 12510
rect 13480 12509 13505 12510
rect 13522 12509 13547 12510
rect 13558 12509 13625 12510
rect 13636 12509 13661 12510
rect 13678 12509 13703 12510
rect 13714 12509 13781 12510
rect 13792 12509 13817 12510
rect 10743 12449 10751 12482
rect 10760 12432 10768 12499
rect 13856 12438 13857 12453
rect 11101 12402 11117 12419
rect 11101 12401 11134 12402
rect 13591 12392 13600 12409
rect 13591 12391 13617 12392
rect 10653 12286 10654 12301
rect 12317 12286 12318 12301
rect 12740 12293 12745 12309
rect 12723 12276 12728 12292
rect 13011 12286 13012 12301
rect 13871 12286 13872 12301
rect 13833 12265 13834 12273
rect 13402 12256 13468 12257
rect 13558 12256 13624 12257
rect 13714 12256 13780 12257
rect 13419 12239 13451 12240
rect 13575 12239 13607 12240
rect 13731 12239 13763 12240
rect 10549 12214 10566 12231
rect 10726 12214 10743 12231
rect 12213 12214 12230 12231
rect 12331 12214 12348 12231
rect 12907 12214 12924 12231
rect 13025 12214 13042 12231
rect 13280 12214 13297 12231
rect 13349 12214 13366 12231
rect 13427 12214 13444 12231
rect 13505 12214 13522 12231
rect 13583 12214 13600 12231
rect 13661 12214 13678 12231
rect 13739 12214 13756 12231
rect 13817 12214 13834 12231
rect 13885 12214 13902 12231
rect 11041 12194 11058 12211
rect 11100 12194 11117 12211
rect 12586 12194 12603 12211
rect 12645 12194 12662 12211
rect 12078 12157 12205 12158
rect 12238 12157 12381 12158
rect 12414 12157 12578 12158
rect 12611 12157 12695 12158
rect 12728 12157 12764 12158
rect 12781 12157 12899 12158
rect 12932 12157 13075 12158
rect 13108 12157 13272 12158
rect 13305 12157 13419 12158
rect 13451 12157 13575 12158
rect 13607 12157 13731 12158
rect 13763 12157 13877 12158
rect 13910 12157 13935 12158
rect 13968 12157 13997 12158
rect 14026 12141 14027 12163
rect 14069 12141 14070 12163
rect 14531 12158 14569 12169
rect 31691 12158 31729 12169
rect 14026 12140 14070 12141
rect 14441 12140 14458 12158
rect 14534 12140 14551 12158
rect 14605 12140 14622 12158
rect 14701 12140 14718 12158
rect 14794 12140 14811 12158
rect 14865 12140 14882 12158
rect 14961 12140 14978 12158
rect 15054 12140 15071 12158
rect 15125 12140 15142 12158
rect 15221 12140 15238 12158
rect 31081 12140 31098 12158
rect 31174 12140 31191 12158
rect 31245 12140 31262 12158
rect 31341 12140 31358 12158
rect 31434 12140 31451 12158
rect 31505 12140 31522 12158
rect 31601 12140 31618 12158
rect 31694 12140 31711 12158
rect 31765 12140 31782 12158
rect 14531 12129 14569 12140
rect 31691 12129 31729 12140
rect 9516 12101 9560 12102
rect 9516 12079 9517 12101
rect 9559 12079 9560 12101
rect 11041 12087 11058 12104
rect 11100 12087 11117 12104
rect 12586 12087 12603 12104
rect 12645 12102 12662 12104
rect 12632 12101 12676 12102
rect 10549 12067 10566 12084
rect 10726 12067 10743 12084
rect 12213 12067 12230 12084
rect 12331 12067 12348 12084
rect 12632 12079 12633 12101
rect 12645 12087 12662 12101
rect 12675 12079 12676 12101
rect 14518 12101 14562 12102
rect 12907 12067 12924 12084
rect 13025 12067 13042 12084
rect 13280 12067 13297 12084
rect 13349 12067 13366 12084
rect 13427 12067 13444 12084
rect 13505 12067 13522 12084
rect 13583 12067 13600 12084
rect 13661 12067 13678 12084
rect 13739 12067 13756 12084
rect 13817 12067 13834 12084
rect 13885 12067 13902 12084
rect 14518 12079 14519 12101
rect 14561 12079 14562 12101
rect 13419 12058 13451 12059
rect 13575 12058 13607 12059
rect 13731 12058 13763 12059
rect 13816 12042 13817 12050
rect 13402 12041 13468 12042
rect 13558 12041 13624 12042
rect 13714 12041 13780 12042
rect 10638 12012 10639 12027
rect 12302 12012 12303 12027
rect 12723 12006 12728 12023
rect 12996 12012 12997 12027
rect 13856 12012 13857 12027
rect 12740 11989 12745 12006
rect 11101 11914 11117 11931
rect 13591 11924 13600 11941
rect 13591 11923 13617 11924
rect 11101 11913 11134 11914
rect 10743 11816 10751 11849
rect 10760 11799 10768 11866
rect 13871 11860 13872 11875
rect 13833 11797 13834 11805
rect 10653 11776 10654 11791
rect 12317 11776 12318 11791
rect 13011 11776 13012 11791
rect 13366 11788 13391 11789
rect 13402 11788 13469 11789
rect 13480 11788 13505 11789
rect 13522 11788 13547 11789
rect 13558 11788 13625 11789
rect 13636 11788 13661 11789
rect 13678 11788 13703 11789
rect 13714 11788 13781 11789
rect 13792 11788 13817 11789
rect 12357 11771 12365 11772
rect 13051 11771 13059 11772
rect 13366 11771 13374 11772
rect 13419 11771 13452 11772
rect 13497 11771 13505 11772
rect 13522 11771 13530 11772
rect 13575 11771 13608 11772
rect 13653 11771 13661 11772
rect 13678 11771 13686 11772
rect 13731 11771 13764 11772
rect 13809 11771 13817 11772
rect 10751 11763 10760 11764
rect 12364 11754 12374 11755
rect 10625 11746 10726 11747
rect 10743 11746 10768 11747
rect 12381 11737 12391 11755
rect 13058 11754 13068 11755
rect 13075 11737 13085 11755
rect 13280 11747 13297 11764
rect 13349 11747 13366 11764
rect 13427 11747 13444 11764
rect 13505 11747 13522 11764
rect 13583 11747 13600 11764
rect 13661 11747 13678 11764
rect 13739 11747 13756 11764
rect 13817 11747 13834 11764
rect 13885 11747 13902 11764
rect 10625 11729 10633 11730
rect 10659 11729 10692 11730
rect 10718 11729 10726 11730
rect 10743 11729 10751 11730
rect 10549 11705 10566 11722
rect 10608 11705 10625 11722
rect 10667 11705 10684 11722
rect 10726 11705 10743 11722
rect 11041 11705 11058 11722
rect 11100 11705 11117 11722
rect 12213 11705 12230 11722
rect 12272 11705 12289 11722
rect 12331 11705 12348 11722
rect 12586 11705 12603 11722
rect 12645 11705 12662 11722
rect 12907 11705 12924 11722
rect 12966 11705 12983 11722
rect 13025 11705 13042 11722
rect 9598 11649 9599 11671
rect 9641 11649 9642 11671
rect 10580 11650 10595 11651
rect 10639 11650 10654 11651
rect 10698 11650 10713 11651
rect 11072 11650 11087 11651
rect 12244 11650 12259 11651
rect 12303 11650 12318 11651
rect 12617 11650 12632 11651
rect 12938 11650 12953 11651
rect 12997 11650 13012 11651
rect 13311 11650 13326 11651
rect 13389 11650 13404 11651
rect 13467 11650 13482 11651
rect 13545 11650 13560 11651
rect 13623 11650 13638 11651
rect 13701 11650 13716 11651
rect 13779 11650 13794 11651
rect 13857 11650 13872 11651
rect 9598 11648 9642 11649
rect 12755 11648 12765 11649
rect 12772 11648 12782 11649
rect 14456 11631 14473 11649
rect 14531 11619 14569 11661
rect 14581 11631 14598 11649
rect 14631 11631 14648 11649
rect 14716 11631 14733 11649
rect 14794 11631 14811 11649
rect 14841 11631 14858 11649
rect 14891 11631 14908 11649
rect 14976 11631 14993 11649
rect 15054 11631 15071 11649
rect 15101 11631 15118 11649
rect 15151 11631 15168 11649
rect 15236 11631 15253 11649
rect 31022 11631 31028 11649
rect 31096 11631 31113 11649
rect 31174 11631 31191 11649
rect 31221 11631 31238 11649
rect 31271 11631 31288 11649
rect 31356 11631 31373 11649
rect 31434 11631 31451 11649
rect 31481 11631 31498 11649
rect 31531 11631 31548 11649
rect 31616 11631 31633 11649
rect 31691 11619 31729 11661
rect 31741 11631 31758 11649
rect 31791 11631 31808 11649
rect 9598 11609 9642 11610
rect 9598 11587 9599 11609
rect 9641 11587 9642 11609
rect 12714 11609 12758 11610
rect 12714 11587 12715 11609
rect 12757 11587 12758 11609
rect 9707 11558 9724 11575
rect 9766 11558 9783 11575
rect 10549 11558 10566 11575
rect 10608 11558 10625 11575
rect 10667 11558 10684 11575
rect 10726 11558 10743 11575
rect 11041 11558 11058 11575
rect 11100 11558 11117 11575
rect 12213 11558 12230 11575
rect 12272 11558 12289 11575
rect 12331 11558 12348 11575
rect 12586 11558 12603 11575
rect 12645 11558 12662 11575
rect 12907 11558 12924 11575
rect 12966 11558 12983 11575
rect 13025 11558 13042 11575
rect 10625 11550 10633 11551
rect 10659 11550 10692 11551
rect 10718 11550 10726 11551
rect 10743 11550 10751 11551
rect 10625 11533 10726 11534
rect 10743 11533 10777 11534
rect 12381 11526 12391 11543
rect 13075 11526 13085 11543
rect 12364 11525 12391 11526
rect 13058 11525 13085 11526
rect 10638 11504 10639 11519
rect 12302 11504 12303 11519
rect 12996 11504 12997 11519
rect 13280 11516 13297 11533
rect 13349 11516 13366 11533
rect 13427 11516 13444 11533
rect 13505 11516 13522 11533
rect 13583 11516 13600 11533
rect 13661 11516 13678 11533
rect 13739 11516 13756 11533
rect 13817 11516 13834 11533
rect 13885 11516 13902 11533
rect 13366 11508 13374 11509
rect 13419 11508 13452 11509
rect 13497 11508 13505 11509
rect 13522 11508 13530 11509
rect 13575 11508 13608 11509
rect 13653 11508 13661 11509
rect 13678 11508 13686 11509
rect 13731 11508 13764 11509
rect 13809 11508 13817 11509
rect 13816 11492 13817 11500
rect 13366 11491 13391 11492
rect 13402 11491 13469 11492
rect 13480 11491 13505 11492
rect 13522 11491 13547 11492
rect 13558 11491 13625 11492
rect 13636 11491 13661 11492
rect 13678 11491 13703 11492
rect 13714 11491 13781 11492
rect 13792 11491 13817 11492
rect 10743 11431 10751 11464
rect 10760 11414 10768 11481
rect 13856 11420 13857 11435
rect 9767 11384 9783 11401
rect 11101 11384 11117 11401
rect 9767 11383 9800 11384
rect 11101 11383 11134 11384
rect 13591 11374 13600 11391
rect 13591 11373 13617 11374
rect 10653 11268 10654 11283
rect 12317 11268 12318 11283
rect 12740 11275 12745 11291
rect 12723 11258 12728 11274
rect 13011 11268 13012 11283
rect 13871 11268 13872 11283
rect 13833 11247 13834 11255
rect 13402 11238 13468 11239
rect 13558 11238 13624 11239
rect 13714 11238 13780 11239
rect 13419 11221 13451 11222
rect 13575 11221 13607 11222
rect 13731 11221 13763 11222
rect 10549 11196 10566 11213
rect 10726 11196 10743 11213
rect 12213 11196 12230 11213
rect 12331 11196 12348 11213
rect 12907 11196 12924 11213
rect 13025 11196 13042 11213
rect 13280 11196 13297 11213
rect 13349 11196 13366 11213
rect 13427 11196 13444 11213
rect 13505 11196 13522 11213
rect 13583 11196 13600 11213
rect 13661 11196 13678 11213
rect 13739 11196 13756 11213
rect 13817 11196 13834 11213
rect 13885 11196 13902 11213
rect 9707 11176 9724 11193
rect 9766 11176 9783 11193
rect 11041 11176 11058 11193
rect 11100 11176 11117 11193
rect 12586 11176 12603 11193
rect 12645 11176 12662 11193
rect 31738 11157 31739 11179
rect 31781 11157 31782 11179
rect 31738 11156 31782 11157
rect 14531 11140 14569 11151
rect 31691 11140 31729 11151
rect 12078 11139 12205 11140
rect 12238 11139 12381 11140
rect 12414 11139 12578 11140
rect 12611 11139 12695 11140
rect 12728 11139 12764 11140
rect 12781 11139 12899 11140
rect 12932 11139 13075 11140
rect 13108 11139 13272 11140
rect 13305 11139 13419 11140
rect 13451 11139 13575 11140
rect 13607 11139 13731 11140
rect 13763 11139 13877 11140
rect 13910 11139 13935 11140
rect 13968 11139 13997 11140
rect 14441 11122 14458 11140
rect 14534 11122 14551 11140
rect 14605 11122 14622 11140
rect 14701 11122 14718 11140
rect 14794 11122 14811 11140
rect 14865 11122 14882 11140
rect 14961 11122 14978 11140
rect 15054 11122 15071 11140
rect 15125 11122 15142 11140
rect 15221 11122 15238 11140
rect 31081 11122 31098 11140
rect 31174 11122 31191 11140
rect 31245 11122 31262 11140
rect 31341 11122 31358 11140
rect 31434 11122 31451 11140
rect 31505 11122 31522 11140
rect 31601 11122 31618 11140
rect 31694 11122 31711 11140
rect 31765 11122 31782 11140
rect 14531 11111 14569 11122
rect 31691 11111 31729 11122
rect 31738 11117 31782 11118
rect 31738 11095 31739 11117
rect 31781 11095 31782 11117
rect 9707 11069 9724 11086
rect 9766 11069 9783 11086
rect 11041 11069 11058 11086
rect 11100 11069 11117 11086
rect 12586 11069 12603 11086
rect 12645 11069 12662 11086
rect 10549 11049 10566 11066
rect 10726 11049 10743 11066
rect 12213 11049 12230 11066
rect 12331 11049 12348 11066
rect 12907 11049 12924 11066
rect 13025 11049 13042 11066
rect 13280 11049 13297 11066
rect 13349 11049 13366 11066
rect 13427 11049 13444 11066
rect 13505 11049 13522 11066
rect 13583 11049 13600 11066
rect 13661 11049 13678 11066
rect 13739 11049 13756 11066
rect 13817 11049 13834 11066
rect 13885 11049 13902 11066
rect 13419 11040 13451 11041
rect 13575 11040 13607 11041
rect 13731 11040 13763 11041
rect 13816 11024 13817 11032
rect 13402 11023 13468 11024
rect 13558 11023 13624 11024
rect 13714 11023 13780 11024
rect 10638 10994 10639 11009
rect 12302 10994 12303 11009
rect 12723 10988 12728 11005
rect 12996 10994 12997 11009
rect 13856 10994 13857 11009
rect 12740 10971 12745 10988
rect 9767 10896 9783 10913
rect 11101 10896 11117 10913
rect 13591 10906 13600 10923
rect 13591 10905 13617 10906
rect 9767 10895 9800 10896
rect 11101 10895 11134 10896
rect 10743 10798 10751 10831
rect 10760 10781 10768 10848
rect 13871 10842 13872 10857
rect 13833 10779 13834 10787
rect 10653 10758 10654 10773
rect 12317 10758 12318 10773
rect 13011 10758 13012 10773
rect 13366 10770 13391 10771
rect 13402 10770 13469 10771
rect 13480 10770 13505 10771
rect 13522 10770 13547 10771
rect 13558 10770 13625 10771
rect 13636 10770 13661 10771
rect 13678 10770 13703 10771
rect 13714 10770 13781 10771
rect 13792 10770 13817 10771
rect 12357 10753 12365 10754
rect 13051 10753 13059 10754
rect 13366 10753 13374 10754
rect 13419 10753 13452 10754
rect 13497 10753 13505 10754
rect 13522 10753 13530 10754
rect 13575 10753 13608 10754
rect 13653 10753 13661 10754
rect 13678 10753 13686 10754
rect 13731 10753 13764 10754
rect 13809 10753 13817 10754
rect 10751 10745 10760 10746
rect 12364 10736 12374 10737
rect 10625 10728 10726 10729
rect 10743 10728 10768 10729
rect 12381 10719 12391 10737
rect 13058 10736 13068 10737
rect 13075 10719 13085 10737
rect 13280 10729 13297 10746
rect 13349 10729 13366 10746
rect 13427 10729 13444 10746
rect 13505 10729 13522 10746
rect 13583 10729 13600 10746
rect 13661 10729 13678 10746
rect 13739 10729 13756 10746
rect 13817 10729 13834 10746
rect 13885 10729 13902 10746
rect 10625 10711 10633 10712
rect 10659 10711 10692 10712
rect 10718 10711 10726 10712
rect 10743 10711 10751 10712
rect 9707 10687 9724 10704
rect 9766 10687 9783 10704
rect 10549 10687 10566 10704
rect 10608 10687 10625 10704
rect 10667 10687 10684 10704
rect 10726 10687 10743 10704
rect 11041 10687 11058 10704
rect 11100 10687 11117 10704
rect 12213 10687 12230 10704
rect 12272 10687 12289 10704
rect 12331 10687 12348 10704
rect 12586 10687 12603 10704
rect 12645 10687 12662 10704
rect 12907 10687 12924 10704
rect 12966 10687 12983 10704
rect 13025 10687 13042 10704
rect 13944 10665 13945 10687
rect 13987 10665 13988 10687
rect 13944 10664 13988 10665
rect 9738 10632 9753 10633
rect 10580 10632 10595 10633
rect 10639 10632 10654 10633
rect 10698 10632 10713 10633
rect 11072 10632 11087 10633
rect 12244 10632 12259 10633
rect 12303 10632 12318 10633
rect 12617 10632 12632 10633
rect 12938 10632 12953 10633
rect 12997 10632 13012 10633
rect 13311 10632 13326 10633
rect 13389 10632 13404 10633
rect 13467 10632 13482 10633
rect 13545 10632 13560 10633
rect 13623 10632 13638 10633
rect 13701 10632 13716 10633
rect 13779 10632 13794 10633
rect 13857 10632 13872 10633
rect 12755 10630 12765 10631
rect 12772 10630 12782 10631
rect 9762 10625 9806 10626
rect 9762 10603 9763 10625
rect 9805 10603 9806 10625
rect 13944 10625 13988 10626
rect 13944 10603 13945 10625
rect 13987 10603 13988 10625
rect 14456 10613 14473 10631
rect 14531 10601 14569 10643
rect 14581 10613 14598 10631
rect 14631 10613 14648 10631
rect 14716 10613 14733 10631
rect 14794 10613 14811 10631
rect 14841 10613 14858 10631
rect 14891 10613 14908 10631
rect 14976 10613 14993 10631
rect 15054 10613 15071 10631
rect 15101 10613 15118 10631
rect 15151 10613 15168 10631
rect 15236 10613 15253 10631
rect 31022 10613 31028 10631
rect 31096 10613 31113 10631
rect 31174 10613 31191 10631
rect 31221 10613 31238 10631
rect 31271 10613 31288 10631
rect 31356 10613 31373 10631
rect 31434 10613 31451 10631
rect 31481 10613 31498 10631
rect 31531 10613 31548 10631
rect 31616 10613 31633 10631
rect 31691 10601 31729 10643
rect 31741 10613 31758 10631
rect 31791 10613 31808 10631
rect 9707 10540 9724 10557
rect 9766 10540 9783 10557
rect 10549 10540 10566 10557
rect 10608 10540 10625 10557
rect 10667 10540 10684 10557
rect 10726 10540 10743 10557
rect 11041 10540 11058 10557
rect 11100 10540 11117 10557
rect 12213 10540 12230 10557
rect 12272 10540 12289 10557
rect 12331 10540 12348 10557
rect 12586 10540 12603 10557
rect 12645 10540 12662 10557
rect 12907 10540 12924 10557
rect 12966 10540 12983 10557
rect 13025 10540 13042 10557
rect 10625 10532 10633 10533
rect 10659 10532 10692 10533
rect 10718 10532 10726 10533
rect 10743 10532 10751 10533
rect 10625 10515 10726 10516
rect 10743 10515 10777 10516
rect 12381 10508 12391 10525
rect 13075 10508 13085 10525
rect 12364 10507 12391 10508
rect 13058 10507 13085 10508
rect 10638 10486 10639 10501
rect 12302 10486 12303 10501
rect 12996 10486 12997 10501
rect 13280 10498 13297 10515
rect 13349 10498 13366 10515
rect 13427 10498 13444 10515
rect 13505 10498 13522 10515
rect 13583 10498 13600 10515
rect 13661 10498 13678 10515
rect 13739 10498 13756 10515
rect 13817 10498 13834 10515
rect 13885 10498 13902 10515
rect 13366 10490 13374 10491
rect 13419 10490 13452 10491
rect 13497 10490 13505 10491
rect 13522 10490 13530 10491
rect 13575 10490 13608 10491
rect 13653 10490 13661 10491
rect 13678 10490 13686 10491
rect 13731 10490 13764 10491
rect 13809 10490 13817 10491
rect 13816 10474 13817 10482
rect 13366 10473 13391 10474
rect 13402 10473 13469 10474
rect 13480 10473 13505 10474
rect 13522 10473 13547 10474
rect 13558 10473 13625 10474
rect 13636 10473 13661 10474
rect 13678 10473 13703 10474
rect 13714 10473 13781 10474
rect 13792 10473 13817 10474
rect 10743 10413 10751 10446
rect 10760 10396 10768 10463
rect 13856 10402 13857 10417
rect 9767 10366 9783 10383
rect 11101 10366 11117 10383
rect 9767 10365 9800 10366
rect 11101 10365 11134 10366
rect 13591 10356 13600 10373
rect 13591 10355 13617 10356
rect 10653 10250 10654 10265
rect 12317 10250 12318 10265
rect 12740 10257 12745 10273
rect 12723 10240 12728 10256
rect 13011 10250 13012 10265
rect 13871 10250 13872 10265
rect 13833 10229 13834 10237
rect 13402 10220 13468 10221
rect 13558 10220 13624 10221
rect 13714 10220 13780 10221
rect 13419 10203 13451 10204
rect 13575 10203 13607 10204
rect 13731 10203 13763 10204
rect 9516 10173 9517 10195
rect 9559 10173 9560 10195
rect 10549 10178 10566 10195
rect 10726 10178 10743 10195
rect 12213 10178 12230 10195
rect 12331 10178 12348 10195
rect 9516 10172 9560 10173
rect 9707 10158 9724 10175
rect 9766 10158 9783 10175
rect 11041 10158 11058 10175
rect 11100 10158 11117 10175
rect 12586 10158 12603 10175
rect 12645 10158 12662 10175
rect 12796 10173 12797 10195
rect 12839 10173 12840 10195
rect 12907 10178 12924 10195
rect 13025 10178 13042 10195
rect 13280 10178 13297 10195
rect 13349 10178 13366 10195
rect 13427 10178 13444 10195
rect 13505 10178 13522 10195
rect 13583 10178 13600 10195
rect 13661 10178 13678 10195
rect 13739 10178 13756 10195
rect 13817 10178 13834 10195
rect 13885 10178 13902 10195
rect 12796 10172 12840 10173
rect 14026 10173 14027 10195
rect 14069 10173 14070 10195
rect 14026 10172 14070 10173
rect 10418 10133 10462 10134
rect 10418 10111 10419 10133
rect 10461 10111 10462 10133
rect 12632 10133 12676 10134
rect 12632 10122 12633 10133
rect 12675 10122 12676 10133
rect 14531 10122 14569 10133
rect 31691 10122 31729 10133
rect 12078 10121 12205 10122
rect 12238 10121 12381 10122
rect 12414 10121 12578 10122
rect 12611 10121 12695 10122
rect 12728 10121 12764 10122
rect 12781 10121 12899 10122
rect 12932 10121 13075 10122
rect 13108 10121 13272 10122
rect 13305 10121 13419 10122
rect 13451 10121 13575 10122
rect 13607 10121 13731 10122
rect 13763 10121 13877 10122
rect 13910 10121 13935 10122
rect 13968 10121 13997 10122
rect 12632 10111 12633 10121
rect 12675 10111 12676 10121
rect 14441 10104 14458 10122
rect 14534 10104 14551 10122
rect 14605 10104 14622 10122
rect 14701 10104 14718 10122
rect 14794 10104 14811 10122
rect 14865 10104 14882 10122
rect 14961 10104 14978 10122
rect 15054 10104 15071 10122
rect 15125 10104 15142 10122
rect 15221 10104 15238 10122
rect 31081 10104 31098 10122
rect 31174 10104 31191 10122
rect 31245 10104 31262 10122
rect 31341 10104 31358 10122
rect 31434 10104 31451 10122
rect 31505 10104 31522 10122
rect 31601 10104 31618 10122
rect 31694 10104 31711 10122
rect 31765 10104 31782 10122
rect 14531 10093 14569 10104
rect 31691 10093 31729 10104
rect 12586 10051 12603 10068
rect 12645 10051 12662 10068
rect 12213 10031 12230 10048
rect 12331 10031 12348 10048
rect 12907 10031 12924 10048
rect 13025 10031 13042 10048
rect 13280 10031 13297 10048
rect 13349 10031 13366 10048
rect 13427 10031 13444 10048
rect 13505 10031 13522 10048
rect 13583 10031 13600 10048
rect 13661 10031 13678 10048
rect 13739 10031 13756 10048
rect 13817 10031 13834 10048
rect 13885 10031 13902 10048
rect 13419 10022 13451 10023
rect 13575 10022 13607 10023
rect 13731 10022 13763 10023
rect 13816 10006 13817 10014
rect 13402 10005 13468 10006
rect 13558 10005 13624 10006
rect 13714 10005 13780 10006
rect 12302 9976 12303 9991
rect 12723 9970 12728 9987
rect 12996 9976 12997 9991
rect 13856 9976 13857 9991
rect 12740 9953 12745 9970
rect 13591 9888 13600 9905
rect 13591 9887 13617 9888
rect 13871 9824 13872 9839
rect 13833 9761 13834 9769
rect 12317 9740 12318 9755
rect 13011 9740 13012 9755
rect 13366 9752 13391 9753
rect 13402 9752 13469 9753
rect 13480 9752 13505 9753
rect 13522 9752 13547 9753
rect 13558 9752 13625 9753
rect 13636 9752 13661 9753
rect 13678 9752 13703 9753
rect 13714 9752 13781 9753
rect 13792 9752 13817 9753
rect 12357 9735 12365 9736
rect 13051 9735 13059 9736
rect 13366 9735 13374 9736
rect 13419 9735 13452 9736
rect 13497 9735 13505 9736
rect 13522 9735 13530 9736
rect 13575 9735 13608 9736
rect 13653 9735 13661 9736
rect 13678 9735 13686 9736
rect 13731 9735 13764 9736
rect 13809 9735 13817 9736
rect 12364 9718 12374 9719
rect 12381 9701 12391 9719
rect 13058 9718 13068 9719
rect 13075 9701 13085 9719
rect 13280 9711 13297 9728
rect 13349 9711 13366 9728
rect 13427 9711 13444 9728
rect 13505 9711 13522 9728
rect 13583 9711 13600 9728
rect 13661 9711 13678 9728
rect 13739 9711 13756 9728
rect 13817 9711 13834 9728
rect 13885 9711 13902 9728
rect 12213 9669 12230 9686
rect 12272 9669 12289 9686
rect 12331 9669 12348 9686
rect 12586 9669 12603 9686
rect 12645 9669 12662 9686
rect 12907 9669 12924 9686
rect 12966 9669 12983 9686
rect 13025 9669 13042 9686
rect 12244 9614 12259 9615
rect 12303 9614 12318 9615
rect 12617 9614 12632 9615
rect 12714 9599 12715 9621
rect 12757 9613 12758 9621
rect 12938 9614 12953 9615
rect 12997 9614 13012 9615
rect 13311 9614 13326 9615
rect 13389 9614 13404 9615
rect 13467 9614 13482 9615
rect 13545 9614 13560 9615
rect 13623 9614 13638 9615
rect 13701 9614 13716 9615
rect 13779 9614 13794 9615
rect 13857 9614 13872 9615
rect 12755 9612 12765 9613
rect 12772 9612 12782 9613
rect 12757 9599 12758 9612
rect 12714 9598 12758 9599
rect 14456 9595 14473 9613
rect 14531 9583 14569 9625
rect 14581 9595 14598 9613
rect 14631 9595 14648 9613
rect 14716 9595 14733 9613
rect 14794 9595 14811 9613
rect 14841 9595 14858 9613
rect 14891 9595 14908 9613
rect 14976 9595 14993 9613
rect 15054 9595 15071 9613
rect 15101 9595 15118 9613
rect 15151 9595 15168 9613
rect 15236 9595 15253 9613
rect 15314 9595 15331 9613
rect 15361 9595 15378 9613
rect 15411 9595 15428 9613
rect 15496 9595 15513 9613
rect 15574 9595 15591 9613
rect 15621 9595 15638 9613
rect 15671 9595 15688 9613
rect 15756 9595 15773 9613
rect 15834 9595 15851 9613
rect 15881 9595 15898 9613
rect 15931 9595 15948 9613
rect 16016 9595 16033 9613
rect 16094 9595 16111 9613
rect 16141 9595 16158 9613
rect 16191 9595 16208 9613
rect 16276 9595 16293 9613
rect 16354 9595 16371 9613
rect 16401 9595 16418 9613
rect 16451 9595 16468 9613
rect 16536 9595 16553 9613
rect 16614 9595 16631 9613
rect 16661 9595 16678 9613
rect 16711 9595 16728 9613
rect 16796 9595 16813 9613
rect 16874 9595 16891 9613
rect 16921 9595 16938 9613
rect 16971 9595 16988 9613
rect 17056 9595 17073 9613
rect 17134 9595 17151 9613
rect 17181 9595 17198 9613
rect 17231 9595 17248 9613
rect 17316 9595 17333 9613
rect 17394 9595 17411 9613
rect 17441 9595 17458 9613
rect 17491 9595 17508 9613
rect 17576 9595 17593 9613
rect 17654 9595 17671 9613
rect 17701 9595 17718 9613
rect 17751 9595 17768 9613
rect 17836 9595 17853 9613
rect 17914 9595 17931 9613
rect 17961 9595 17978 9613
rect 18011 9595 18028 9613
rect 18096 9595 18113 9613
rect 18174 9595 18191 9613
rect 18221 9595 18238 9613
rect 18271 9595 18288 9613
rect 18356 9595 18373 9613
rect 18434 9595 18451 9613
rect 18481 9595 18498 9613
rect 18531 9595 18548 9613
rect 18616 9595 18633 9613
rect 18694 9595 18711 9613
rect 18741 9595 18758 9613
rect 18791 9595 18808 9613
rect 18876 9595 18893 9613
rect 18954 9595 18971 9613
rect 19001 9595 19018 9613
rect 19051 9595 19068 9613
rect 19136 9595 19153 9613
rect 19214 9595 19231 9613
rect 19261 9595 19278 9613
rect 19311 9595 19328 9613
rect 19396 9595 19413 9613
rect 19474 9595 19491 9613
rect 19521 9595 19538 9613
rect 19571 9595 19588 9613
rect 19656 9595 19673 9613
rect 19734 9595 19751 9613
rect 19781 9595 19798 9613
rect 19831 9595 19848 9613
rect 19916 9595 19933 9613
rect 19994 9595 20011 9613
rect 20041 9595 20058 9613
rect 20091 9595 20108 9613
rect 30240 9595 30248 9613
rect 30316 9595 30333 9613
rect 30394 9595 30411 9613
rect 30441 9595 30458 9613
rect 30491 9595 30508 9613
rect 30576 9595 30593 9613
rect 30654 9595 30671 9613
rect 30701 9595 30718 9613
rect 30751 9595 30768 9613
rect 30836 9595 30853 9613
rect 30914 9595 30931 9613
rect 30961 9595 30978 9613
rect 31011 9595 31028 9613
rect 31096 9595 31113 9613
rect 31174 9595 31191 9613
rect 31221 9595 31238 9613
rect 31271 9595 31288 9613
rect 31356 9595 31373 9613
rect 31434 9595 31451 9613
rect 31481 9595 31498 9613
rect 31531 9595 31548 9613
rect 31616 9595 31633 9613
rect 31691 9583 31729 9625
rect 31741 9595 31758 9613
rect 31791 9595 31808 9613
rect 12796 9559 12840 9560
rect 12213 9522 12230 9539
rect 12272 9522 12289 9539
rect 12331 9522 12348 9539
rect 12586 9522 12603 9539
rect 12645 9522 12662 9539
rect 12796 9537 12797 9559
rect 12839 9537 12840 9559
rect 12907 9522 12924 9539
rect 12966 9522 12983 9539
rect 13025 9522 13042 9539
rect 12381 9490 12391 9507
rect 13075 9490 13085 9507
rect 12364 9489 12391 9490
rect 13058 9489 13085 9490
rect 12302 9468 12303 9483
rect 12996 9468 12997 9483
rect 13280 9480 13297 9497
rect 13349 9480 13366 9497
rect 13427 9480 13444 9497
rect 13505 9480 13522 9497
rect 13583 9480 13600 9497
rect 13661 9480 13678 9497
rect 13739 9480 13756 9497
rect 13817 9480 13834 9497
rect 13885 9480 13902 9497
rect 13366 9472 13374 9473
rect 13419 9472 13452 9473
rect 13497 9472 13505 9473
rect 13522 9472 13530 9473
rect 13575 9472 13608 9473
rect 13653 9472 13661 9473
rect 13678 9472 13686 9473
rect 13731 9472 13764 9473
rect 13809 9472 13817 9473
rect 13816 9456 13817 9464
rect 13366 9455 13391 9456
rect 13402 9455 13469 9456
rect 13480 9455 13505 9456
rect 13522 9455 13547 9456
rect 13558 9455 13625 9456
rect 13636 9455 13661 9456
rect 13678 9455 13703 9456
rect 13714 9455 13781 9456
rect 13792 9455 13817 9456
rect 13856 9384 13857 9399
rect 13591 9338 13600 9355
rect 13591 9337 13617 9338
rect 12317 9232 12318 9247
rect 12740 9239 12745 9255
rect 12723 9222 12728 9238
rect 13011 9232 13012 9247
rect 13871 9232 13872 9247
rect 13833 9211 13834 9219
rect 13402 9202 13468 9203
rect 13558 9202 13624 9203
rect 13714 9202 13780 9203
rect 13419 9185 13451 9186
rect 13575 9185 13607 9186
rect 13731 9185 13763 9186
rect 12213 9160 12230 9177
rect 12331 9160 12348 9177
rect 12907 9160 12924 9177
rect 13025 9160 13042 9177
rect 13280 9160 13297 9177
rect 13349 9160 13366 9177
rect 13427 9160 13444 9177
rect 13505 9160 13522 9177
rect 13583 9160 13600 9177
rect 13661 9160 13678 9177
rect 13739 9160 13756 9177
rect 13817 9160 13834 9177
rect 13885 9160 13902 9177
rect 12586 9140 12603 9157
rect 12645 9140 12662 9157
rect 14531 9104 14569 9115
rect 31691 9104 31729 9115
rect 12078 9103 12205 9104
rect 12238 9103 12381 9104
rect 12414 9103 12578 9104
rect 12611 9103 12695 9104
rect 12728 9103 12764 9104
rect 12781 9103 12899 9104
rect 12932 9103 13075 9104
rect 13108 9103 13272 9104
rect 13305 9103 13419 9104
rect 13451 9103 13575 9104
rect 13607 9103 13731 9104
rect 13763 9103 13877 9104
rect 13910 9103 13935 9104
rect 13968 9103 13997 9104
rect 14441 9086 14458 9104
rect 14534 9086 14551 9104
rect 14605 9086 14622 9104
rect 14701 9086 14718 9104
rect 14794 9086 14811 9104
rect 14865 9086 14882 9104
rect 14961 9086 14978 9104
rect 15054 9086 15071 9104
rect 15125 9086 15142 9104
rect 15221 9086 15238 9104
rect 15314 9086 15331 9104
rect 15385 9086 15402 9104
rect 15481 9086 15498 9104
rect 15574 9086 15591 9104
rect 15645 9086 15662 9104
rect 15741 9086 15758 9104
rect 15834 9086 15851 9104
rect 15905 9086 15922 9104
rect 16001 9086 16018 9104
rect 16094 9086 16111 9104
rect 16165 9086 16182 9104
rect 16261 9086 16278 9104
rect 16354 9086 16371 9104
rect 16425 9086 16442 9104
rect 16521 9086 16538 9104
rect 16614 9086 16631 9104
rect 16685 9086 16702 9104
rect 16781 9086 16798 9104
rect 16874 9086 16891 9104
rect 16945 9086 16962 9104
rect 17041 9086 17058 9104
rect 17134 9086 17151 9104
rect 17205 9086 17222 9104
rect 17301 9086 17318 9104
rect 17394 9086 17411 9104
rect 17465 9086 17482 9104
rect 17561 9086 17578 9104
rect 17654 9086 17671 9104
rect 17725 9086 17742 9104
rect 17821 9086 17838 9104
rect 17914 9086 17931 9104
rect 17985 9086 18002 9104
rect 18081 9086 18098 9104
rect 18174 9086 18191 9104
rect 18245 9086 18262 9104
rect 18341 9086 18358 9104
rect 18434 9086 18451 9104
rect 18505 9086 18522 9104
rect 18601 9086 18618 9104
rect 18694 9086 18711 9104
rect 18765 9086 18782 9104
rect 18861 9086 18878 9104
rect 18954 9086 18971 9104
rect 19025 9086 19042 9104
rect 19121 9086 19138 9104
rect 19214 9086 19231 9104
rect 19285 9086 19302 9104
rect 19381 9086 19398 9104
rect 19474 9086 19491 9104
rect 19545 9086 19562 9104
rect 19641 9086 19658 9104
rect 19734 9086 19751 9104
rect 19805 9086 19822 9104
rect 19901 9086 19918 9104
rect 19994 9086 20011 9104
rect 20065 9086 20082 9104
rect 30301 9086 30318 9104
rect 30394 9086 30411 9104
rect 30465 9086 30482 9104
rect 30561 9086 30578 9104
rect 30654 9086 30671 9104
rect 30725 9086 30742 9104
rect 30821 9086 30838 9104
rect 30914 9086 30931 9104
rect 30985 9086 31002 9104
rect 31081 9086 31098 9104
rect 31174 9086 31191 9104
rect 31245 9086 31262 9104
rect 31341 9086 31358 9104
rect 31434 9086 31451 9104
rect 31505 9086 31522 9104
rect 31601 9086 31618 9104
rect 31694 9086 31711 9104
rect 31765 9086 31782 9104
rect 14531 9075 14569 9086
rect 31691 9075 31729 9086
rect 9844 9067 9888 9068
rect 9844 9045 9845 9067
rect 9887 9045 9888 9067
rect 31656 9067 31700 9068
rect 11041 9033 11058 9050
rect 11100 9033 11117 9050
rect 12586 9033 12603 9050
rect 12645 9033 12662 9050
rect 31656 9045 31657 9067
rect 31699 9045 31700 9067
rect 10668 9013 10685 9030
rect 10786 9013 10803 9030
rect 12213 9013 12230 9030
rect 12331 9013 12348 9030
rect 12907 9013 12924 9030
rect 13025 9013 13042 9030
rect 13280 9013 13297 9030
rect 13349 9013 13366 9030
rect 13427 9013 13444 9030
rect 13505 9013 13522 9030
rect 13583 9013 13600 9030
rect 13661 9013 13678 9030
rect 13739 9013 13756 9030
rect 13817 9013 13834 9030
rect 13885 9013 13902 9030
rect 13419 9004 13451 9005
rect 13575 9004 13607 9005
rect 13731 9004 13763 9005
rect 13816 8988 13817 8996
rect 13402 8987 13468 8988
rect 13558 8987 13624 8988
rect 13714 8987 13780 8988
rect 10757 8958 10758 8973
rect 12302 8958 12303 8973
rect 12723 8952 12728 8969
rect 12996 8958 12997 8973
rect 13856 8958 13857 8973
rect 12740 8935 12745 8952
rect 11101 8860 11117 8877
rect 13591 8870 13600 8887
rect 13591 8869 13617 8870
rect 11101 8859 11134 8860
rect 13871 8806 13872 8821
rect 13833 8743 13834 8751
rect 10772 8722 10773 8737
rect 12317 8722 12318 8737
rect 13011 8722 13012 8737
rect 13366 8734 13391 8735
rect 13402 8734 13469 8735
rect 13480 8734 13505 8735
rect 13522 8734 13547 8735
rect 13558 8734 13625 8735
rect 13636 8734 13661 8735
rect 13678 8734 13703 8735
rect 13714 8734 13781 8735
rect 13792 8734 13817 8735
rect 10812 8717 10820 8718
rect 12357 8717 12365 8718
rect 13051 8717 13059 8718
rect 13366 8717 13374 8718
rect 13419 8717 13452 8718
rect 13497 8717 13505 8718
rect 13522 8717 13530 8718
rect 13575 8717 13608 8718
rect 13653 8717 13661 8718
rect 13678 8717 13686 8718
rect 13731 8717 13764 8718
rect 13809 8717 13817 8718
rect 10819 8700 10829 8701
rect 10836 8683 10846 8701
rect 12364 8700 12374 8701
rect 12381 8683 12391 8701
rect 13058 8700 13068 8701
rect 13075 8683 13085 8701
rect 13280 8693 13297 8710
rect 13349 8693 13366 8710
rect 13427 8693 13444 8710
rect 13505 8693 13522 8710
rect 13583 8693 13600 8710
rect 13661 8693 13678 8710
rect 13739 8693 13756 8710
rect 13817 8693 13834 8710
rect 13885 8693 13902 8710
rect 10668 8651 10685 8668
rect 10727 8651 10744 8668
rect 10786 8651 10803 8668
rect 11041 8651 11058 8668
rect 11100 8651 11117 8668
rect 12213 8651 12230 8668
rect 12272 8651 12289 8668
rect 12331 8651 12348 8668
rect 12586 8651 12603 8668
rect 12645 8651 12662 8668
rect 12907 8651 12924 8668
rect 12966 8651 12983 8668
rect 13025 8651 13042 8668
rect 13944 8615 13945 8637
rect 13987 8615 13988 8637
rect 13944 8614 13988 8615
rect 10699 8596 10714 8597
rect 10758 8596 10773 8597
rect 11072 8596 11087 8597
rect 12244 8596 12259 8597
rect 12303 8596 12318 8597
rect 12617 8596 12632 8597
rect 12938 8596 12953 8597
rect 12997 8596 13012 8597
rect 13311 8596 13326 8597
rect 13389 8596 13404 8597
rect 13467 8596 13482 8597
rect 13545 8596 13560 8597
rect 13623 8596 13638 8597
rect 13701 8596 13716 8597
rect 13779 8596 13794 8597
rect 13857 8596 13872 8597
rect 12755 8594 12765 8595
rect 12772 8594 12782 8595
rect 14456 8577 14473 8595
rect 9762 8575 9806 8576
rect 9762 8553 9763 8575
rect 9805 8553 9806 8575
rect 12714 8575 12758 8576
rect 12714 8553 12715 8575
rect 12757 8553 12758 8575
rect 14026 8575 14070 8576
rect 14026 8553 14027 8575
rect 14069 8553 14070 8575
rect 14531 8565 14569 8607
rect 14581 8577 14598 8595
rect 14631 8577 14648 8595
rect 14716 8577 14733 8595
rect 14794 8577 14811 8595
rect 14841 8577 14858 8595
rect 14891 8577 14908 8595
rect 14976 8577 14993 8595
rect 15054 8577 15071 8595
rect 15101 8577 15118 8595
rect 15151 8577 15168 8595
rect 15236 8577 15253 8595
rect 15314 8577 15331 8595
rect 15361 8577 15378 8595
rect 15411 8577 15428 8595
rect 15496 8577 15513 8595
rect 15574 8577 15591 8595
rect 15621 8577 15638 8595
rect 15671 8577 15688 8595
rect 15756 8577 15773 8595
rect 15834 8577 15851 8595
rect 15881 8577 15898 8595
rect 15931 8577 15948 8595
rect 16016 8577 16033 8595
rect 16094 8577 16111 8595
rect 16141 8577 16158 8595
rect 16191 8577 16208 8595
rect 16276 8577 16293 8595
rect 16354 8577 16371 8595
rect 16401 8577 16418 8595
rect 16451 8577 16468 8595
rect 16536 8577 16553 8595
rect 16614 8577 16631 8595
rect 16661 8577 16678 8595
rect 16711 8577 16728 8595
rect 16796 8577 16813 8595
rect 16874 8577 16891 8595
rect 16921 8577 16938 8595
rect 16971 8577 16988 8595
rect 17056 8577 17073 8595
rect 17134 8577 17151 8595
rect 17181 8577 17198 8595
rect 17231 8577 17248 8595
rect 17316 8577 17333 8595
rect 17394 8577 17411 8595
rect 17441 8577 17458 8595
rect 17491 8577 17508 8595
rect 17576 8577 17593 8595
rect 17654 8577 17671 8595
rect 17701 8577 17718 8595
rect 17751 8577 17768 8595
rect 17836 8577 17853 8595
rect 17914 8577 17931 8595
rect 17961 8577 17978 8595
rect 18011 8577 18028 8595
rect 18096 8577 18113 8595
rect 18174 8577 18191 8595
rect 18221 8577 18238 8595
rect 18271 8577 18288 8595
rect 18356 8577 18373 8595
rect 18434 8577 18451 8595
rect 18481 8577 18498 8595
rect 18531 8577 18548 8595
rect 18616 8577 18633 8595
rect 18694 8577 18711 8595
rect 18741 8577 18758 8595
rect 18791 8577 18808 8595
rect 18876 8577 18893 8595
rect 18954 8577 18971 8595
rect 19001 8577 19018 8595
rect 19051 8577 19068 8595
rect 19136 8577 19153 8595
rect 19214 8577 19231 8595
rect 19261 8577 19278 8595
rect 19311 8577 19328 8595
rect 19396 8577 19413 8595
rect 19474 8577 19491 8595
rect 19521 8577 19538 8595
rect 19571 8577 19588 8595
rect 19656 8577 19673 8595
rect 19734 8577 19751 8595
rect 19781 8577 19798 8595
rect 19831 8577 19848 8595
rect 19916 8577 19933 8595
rect 19994 8577 20011 8595
rect 20041 8577 20058 8595
rect 20091 8577 20108 8595
rect 30240 8577 30248 8595
rect 30316 8577 30333 8595
rect 30394 8577 30411 8595
rect 30441 8577 30458 8595
rect 30491 8577 30508 8595
rect 30576 8577 30593 8595
rect 30654 8577 30671 8595
rect 30701 8577 30718 8595
rect 30751 8577 30768 8595
rect 30836 8577 30853 8595
rect 30914 8577 30931 8595
rect 30961 8577 30978 8595
rect 31011 8577 31028 8595
rect 31096 8577 31113 8595
rect 31174 8577 31191 8595
rect 31221 8577 31238 8595
rect 31271 8577 31288 8595
rect 31356 8577 31373 8595
rect 31434 8577 31451 8595
rect 31481 8577 31498 8595
rect 31531 8577 31548 8595
rect 31616 8577 31633 8595
rect 31691 8565 31729 8607
rect 31741 8577 31758 8595
rect 31791 8577 31808 8595
rect 10668 8504 10685 8521
rect 10727 8504 10744 8521
rect 10786 8504 10803 8521
rect 11041 8504 11058 8521
rect 11100 8504 11117 8521
rect 12213 8504 12230 8521
rect 12272 8504 12289 8521
rect 12331 8504 12348 8521
rect 12586 8504 12603 8521
rect 12645 8504 12662 8521
rect 12907 8504 12924 8521
rect 12966 8504 12983 8521
rect 13025 8504 13042 8521
rect 10836 8472 10846 8489
rect 12381 8472 12391 8489
rect 13075 8472 13085 8489
rect 10819 8471 10846 8472
rect 12364 8471 12391 8472
rect 13058 8471 13085 8472
rect 10757 8450 10758 8465
rect 12302 8450 12303 8465
rect 12996 8450 12997 8465
rect 13280 8462 13297 8479
rect 13349 8462 13366 8479
rect 13427 8462 13444 8479
rect 13505 8462 13522 8479
rect 13583 8462 13600 8479
rect 13661 8462 13678 8479
rect 13739 8462 13756 8479
rect 13817 8462 13834 8479
rect 13885 8462 13902 8479
rect 13366 8454 13374 8455
rect 13419 8454 13452 8455
rect 13497 8454 13505 8455
rect 13522 8454 13530 8455
rect 13575 8454 13608 8455
rect 13653 8454 13661 8455
rect 13678 8454 13686 8455
rect 13731 8454 13764 8455
rect 13809 8454 13817 8455
rect 13816 8438 13817 8446
rect 13366 8437 13391 8438
rect 13402 8437 13469 8438
rect 13480 8437 13505 8438
rect 13522 8437 13547 8438
rect 13558 8437 13625 8438
rect 13636 8437 13661 8438
rect 13678 8437 13703 8438
rect 13714 8437 13781 8438
rect 13792 8437 13817 8438
rect 13856 8366 13857 8381
rect 11101 8330 11117 8347
rect 11101 8329 11134 8330
rect 13591 8320 13600 8337
rect 13591 8319 13617 8320
rect 10772 8214 10773 8229
rect 12317 8214 12318 8229
rect 12740 8221 12745 8237
rect 12723 8204 12728 8220
rect 13011 8214 13012 8229
rect 13871 8214 13872 8229
rect 13833 8193 13834 8201
rect 13402 8184 13468 8185
rect 13558 8184 13624 8185
rect 13714 8184 13780 8185
rect 13419 8167 13451 8168
rect 13575 8167 13607 8168
rect 13731 8167 13763 8168
rect 10668 8142 10685 8159
rect 10786 8142 10803 8159
rect 12213 8142 12230 8159
rect 12331 8142 12348 8159
rect 11041 8122 11058 8139
rect 11100 8122 11117 8139
rect 12586 8122 12603 8139
rect 12632 8123 12633 8145
rect 12645 8123 12662 8139
rect 12675 8123 12676 8145
rect 12907 8142 12924 8159
rect 13025 8142 13042 8159
rect 13280 8142 13297 8159
rect 13349 8142 13366 8159
rect 13427 8142 13444 8159
rect 13505 8142 13522 8159
rect 13583 8142 13600 8159
rect 13661 8142 13678 8159
rect 13739 8142 13756 8159
rect 13817 8142 13834 8159
rect 12632 8122 12676 8123
rect 13862 8123 13863 8145
rect 13885 8142 13902 8159
rect 13905 8123 13906 8145
rect 13862 8122 13906 8123
rect 14531 8086 14569 8097
rect 31691 8086 31729 8097
rect 12078 8085 12205 8086
rect 12238 8085 12381 8086
rect 12414 8085 12578 8086
rect 12611 8085 12695 8086
rect 12728 8085 12764 8086
rect 12781 8085 12899 8086
rect 12932 8085 13075 8086
rect 13108 8085 13272 8086
rect 13305 8085 13419 8086
rect 13451 8085 13575 8086
rect 13607 8085 13731 8086
rect 13763 8085 13877 8086
rect 13910 8085 13935 8086
rect 13968 8085 13997 8086
rect 9844 8083 9888 8084
rect 9844 8061 9845 8083
rect 9887 8061 9888 8083
rect 12632 8083 12676 8084
rect 12632 8061 12633 8083
rect 12675 8061 12676 8083
rect 14441 8068 14458 8086
rect 14534 8068 14551 8086
rect 14605 8068 14622 8086
rect 14701 8068 14718 8086
rect 14794 8068 14811 8086
rect 14865 8068 14882 8086
rect 14961 8068 14978 8086
rect 15054 8068 15071 8086
rect 15125 8068 15142 8086
rect 15221 8068 15238 8086
rect 15314 8068 15331 8086
rect 15385 8068 15402 8086
rect 15481 8068 15498 8086
rect 15574 8068 15591 8086
rect 15645 8068 15662 8086
rect 15741 8068 15758 8086
rect 15834 8068 15851 8086
rect 15905 8068 15922 8086
rect 16001 8068 16018 8086
rect 16094 8068 16111 8086
rect 16165 8068 16182 8086
rect 16261 8068 16278 8086
rect 16354 8068 16371 8086
rect 16425 8068 16442 8086
rect 16521 8068 16538 8086
rect 16614 8068 16631 8086
rect 16685 8068 16702 8086
rect 16781 8068 16798 8086
rect 16874 8068 16891 8086
rect 16945 8068 16962 8086
rect 17041 8068 17058 8086
rect 17134 8068 17151 8086
rect 17205 8068 17222 8086
rect 17301 8068 17318 8086
rect 17394 8068 17411 8086
rect 17465 8068 17482 8086
rect 17561 8068 17578 8086
rect 17654 8068 17671 8086
rect 17725 8068 17742 8086
rect 17821 8068 17838 8086
rect 17914 8068 17931 8086
rect 17985 8068 18002 8086
rect 18081 8068 18098 8086
rect 18174 8068 18191 8086
rect 18245 8068 18262 8086
rect 18341 8068 18358 8086
rect 18434 8068 18451 8086
rect 18505 8068 18522 8086
rect 18601 8068 18618 8086
rect 18694 8068 18711 8086
rect 18765 8068 18782 8086
rect 18861 8068 18878 8086
rect 18954 8068 18971 8086
rect 19025 8068 19042 8086
rect 19121 8068 19138 8086
rect 19214 8068 19231 8086
rect 19285 8068 19302 8086
rect 19381 8068 19398 8086
rect 19474 8068 19491 8086
rect 19545 8068 19562 8086
rect 19641 8068 19658 8086
rect 19734 8068 19751 8086
rect 19805 8068 19822 8086
rect 19901 8068 19918 8086
rect 19994 8068 20011 8086
rect 20065 8068 20082 8086
rect 30301 8068 30318 8086
rect 30394 8068 30411 8086
rect 30465 8068 30482 8086
rect 30561 8068 30578 8086
rect 30654 8068 30671 8086
rect 30725 8068 30742 8086
rect 30821 8068 30838 8086
rect 30914 8068 30931 8086
rect 30985 8068 31002 8086
rect 31081 8068 31098 8086
rect 31174 8068 31191 8086
rect 31245 8068 31262 8086
rect 31341 8068 31358 8086
rect 31434 8068 31451 8086
rect 31505 8068 31522 8086
rect 31601 8068 31618 8086
rect 31694 8068 31711 8086
rect 31765 8068 31782 8086
rect 14531 8057 14569 8068
rect 31691 8057 31729 8068
rect 9958 8015 9975 8032
rect 10017 8015 10034 8032
rect 11041 8015 11058 8032
rect 11100 8015 11117 8032
rect 12586 8015 12603 8032
rect 12645 8015 12662 8032
rect 1146 7997 2716 7998
rect 10668 7995 10685 8012
rect 10786 7995 10803 8012
rect 12213 7995 12230 8012
rect 12331 7995 12348 8012
rect 12907 7995 12924 8012
rect 13025 7995 13042 8012
rect 13280 7995 13297 8012
rect 13349 7995 13366 8012
rect 13427 7995 13444 8012
rect 13505 7995 13522 8012
rect 13583 7995 13600 8012
rect 13661 7995 13678 8012
rect 13739 7995 13756 8012
rect 13817 7995 13834 8012
rect 13885 7995 13902 8012
rect 13419 7986 13451 7987
rect 13575 7986 13607 7987
rect 13731 7986 13763 7987
rect 13816 7970 13817 7978
rect 13402 7969 13468 7970
rect 13558 7969 13624 7970
rect 13714 7969 13780 7970
rect 1281 7927 1298 7944
rect 1340 7927 1357 7944
rect 1595 7927 1612 7944
rect 1654 7927 1671 7944
rect 1909 7927 1926 7944
rect 1968 7927 1985 7944
rect 2223 7927 2240 7944
rect 2282 7927 2299 7944
rect 2537 7927 2554 7944
rect 2596 7927 2613 7944
rect 10757 7940 10758 7955
rect 12302 7940 12303 7955
rect 12723 7934 12728 7951
rect 12996 7940 12997 7955
rect 13856 7940 13857 7955
rect 12740 7917 12745 7934
rect 1379 7835 1434 7844
rect 1579 7826 1675 7844
rect 1693 7835 1748 7844
rect 1893 7826 1989 7844
rect 2007 7835 2062 7844
rect 2207 7826 2303 7844
rect 2321 7835 2376 7844
rect 2521 7826 2617 7844
rect 2635 7835 2690 7844
rect 10018 7842 10034 7859
rect 11101 7842 11117 7859
rect 13591 7852 13600 7869
rect 13591 7851 13617 7852
rect 10018 7841 10051 7842
rect 11101 7841 11134 7842
rect 1179 7818 1223 7819
rect 1179 7776 1180 7818
rect 1222 7776 1223 7818
rect 1357 7805 1366 7806
rect 1671 7805 1680 7806
rect 1985 7805 1994 7806
rect 2299 7805 2308 7806
rect 2613 7805 2622 7806
rect 13871 7788 13872 7803
rect 1179 7775 1187 7776
rect 1215 7775 1223 7776
rect 13833 7725 13834 7733
rect 10772 7704 10773 7719
rect 12317 7704 12318 7719
rect 13011 7704 13012 7719
rect 13366 7716 13391 7717
rect 13402 7716 13469 7717
rect 13480 7716 13505 7717
rect 13522 7716 13547 7717
rect 13558 7716 13625 7717
rect 13636 7716 13661 7717
rect 13678 7716 13703 7717
rect 13714 7716 13781 7717
rect 13792 7716 13817 7717
rect 10812 7699 10820 7700
rect 12357 7699 12365 7700
rect 13051 7699 13059 7700
rect 13366 7699 13374 7700
rect 13419 7699 13452 7700
rect 13497 7699 13505 7700
rect 13522 7699 13530 7700
rect 13575 7699 13608 7700
rect 13653 7699 13661 7700
rect 13678 7699 13686 7700
rect 13731 7699 13764 7700
rect 13809 7699 13817 7700
rect 10819 7682 10829 7683
rect 1281 7649 1298 7666
rect 1340 7649 1357 7666
rect 1595 7649 1612 7666
rect 1654 7649 1671 7666
rect 1909 7649 1926 7666
rect 1968 7649 1985 7666
rect 2223 7649 2240 7666
rect 2282 7649 2299 7666
rect 2537 7649 2554 7666
rect 2596 7649 2613 7666
rect 10836 7665 10846 7683
rect 12364 7682 12374 7683
rect 12381 7665 12391 7683
rect 13058 7682 13068 7683
rect 13075 7665 13085 7683
rect 13280 7675 13297 7692
rect 13349 7675 13366 7692
rect 13427 7675 13444 7692
rect 13505 7675 13522 7692
rect 13583 7675 13600 7692
rect 13661 7675 13678 7692
rect 13739 7675 13756 7692
rect 13817 7675 13834 7692
rect 13885 7675 13902 7692
rect 9958 7633 9975 7650
rect 10017 7633 10034 7650
rect 10668 7633 10685 7650
rect 10727 7633 10744 7650
rect 10786 7633 10803 7650
rect 11041 7633 11058 7650
rect 11100 7633 11117 7650
rect 12213 7633 12230 7650
rect 12272 7633 12289 7650
rect 12331 7633 12348 7650
rect 12586 7633 12603 7650
rect 12645 7633 12662 7650
rect 12907 7633 12924 7650
rect 12966 7633 12983 7650
rect 13025 7633 13042 7650
rect 1146 7591 1273 7592
rect 1306 7591 1390 7592
rect 1423 7591 1587 7592
rect 1620 7591 1704 7592
rect 1737 7591 1901 7592
rect 1934 7591 2018 7592
rect 2051 7591 2215 7592
rect 2248 7591 2332 7592
rect 2365 7591 2529 7592
rect 2562 7591 2646 7592
rect 2679 7591 2716 7592
rect 9989 7578 10004 7579
rect 10699 7578 10714 7579
rect 10758 7578 10773 7579
rect 11072 7578 11087 7579
rect 12244 7578 12259 7579
rect 12303 7578 12318 7579
rect 12617 7578 12632 7579
rect 12938 7578 12953 7579
rect 12997 7578 13012 7579
rect 13311 7578 13326 7579
rect 13389 7578 13404 7579
rect 13467 7578 13482 7579
rect 13545 7578 13560 7579
rect 13623 7578 13638 7579
rect 13701 7578 13716 7579
rect 13779 7578 13794 7579
rect 13857 7578 13872 7579
rect 12755 7576 12765 7577
rect 12772 7576 12782 7577
rect 14456 7559 14473 7577
rect 14531 7547 14569 7589
rect 14581 7559 14598 7577
rect 14631 7559 14648 7577
rect 14716 7559 14733 7577
rect 14794 7559 14811 7577
rect 14841 7559 14858 7577
rect 14891 7559 14908 7577
rect 14976 7559 14993 7577
rect 15054 7559 15071 7577
rect 15101 7559 15118 7577
rect 15151 7559 15168 7577
rect 15236 7559 15253 7577
rect 15314 7559 15331 7577
rect 15361 7559 15378 7577
rect 15411 7559 15428 7577
rect 15496 7559 15513 7577
rect 15574 7559 15591 7577
rect 15621 7559 15638 7577
rect 15671 7559 15688 7577
rect 15756 7559 15773 7577
rect 15834 7559 15851 7577
rect 15881 7559 15898 7577
rect 15931 7559 15948 7577
rect 16016 7559 16033 7577
rect 16094 7559 16111 7577
rect 16141 7559 16158 7577
rect 16191 7559 16208 7577
rect 16276 7559 16293 7577
rect 16354 7559 16371 7577
rect 16401 7559 16418 7577
rect 16451 7559 16468 7577
rect 16536 7559 16553 7577
rect 16614 7559 16631 7577
rect 16661 7559 16678 7577
rect 16711 7559 16728 7577
rect 16796 7559 16813 7577
rect 16874 7559 16891 7577
rect 16921 7559 16938 7577
rect 16971 7559 16988 7577
rect 17056 7559 17073 7577
rect 17134 7559 17151 7577
rect 17181 7559 17198 7577
rect 17231 7559 17248 7577
rect 17316 7559 17333 7577
rect 17394 7559 17411 7577
rect 17441 7559 17458 7577
rect 17491 7559 17508 7577
rect 17576 7559 17593 7577
rect 17654 7559 17671 7577
rect 17701 7559 17718 7577
rect 17751 7559 17768 7577
rect 17836 7559 17853 7577
rect 17914 7559 17931 7577
rect 17961 7559 17978 7577
rect 18011 7559 18028 7577
rect 18096 7559 18113 7577
rect 18174 7559 18191 7577
rect 18221 7559 18238 7577
rect 18271 7559 18288 7577
rect 18356 7559 18373 7577
rect 18434 7559 18451 7577
rect 18481 7559 18498 7577
rect 18531 7559 18548 7577
rect 18616 7559 18633 7577
rect 18694 7559 18711 7577
rect 18741 7559 18758 7577
rect 18791 7559 18808 7577
rect 18876 7559 18893 7577
rect 18954 7559 18971 7577
rect 19001 7559 19018 7577
rect 19051 7559 19068 7577
rect 19136 7559 19153 7577
rect 19214 7559 19231 7577
rect 19261 7559 19278 7577
rect 19311 7559 19328 7577
rect 19396 7559 19413 7577
rect 19474 7559 19491 7577
rect 19521 7559 19538 7577
rect 19571 7559 19588 7577
rect 19656 7559 19673 7577
rect 19734 7559 19751 7577
rect 19781 7559 19798 7577
rect 19831 7559 19848 7577
rect 19916 7559 19933 7577
rect 19994 7559 20011 7577
rect 20041 7559 20058 7577
rect 20091 7559 20108 7577
rect 30240 7559 30248 7577
rect 30316 7559 30333 7577
rect 30394 7559 30411 7577
rect 30441 7559 30458 7577
rect 30491 7559 30508 7577
rect 30576 7559 30593 7577
rect 30654 7559 30671 7577
rect 30701 7559 30718 7577
rect 30751 7559 30768 7577
rect 30836 7559 30853 7577
rect 30914 7559 30931 7577
rect 30961 7559 30978 7577
rect 31011 7559 31028 7577
rect 31096 7559 31113 7577
rect 31174 7559 31191 7577
rect 31221 7559 31238 7577
rect 31271 7559 31288 7577
rect 31356 7559 31373 7577
rect 31434 7559 31451 7577
rect 31481 7559 31498 7577
rect 31531 7559 31548 7577
rect 31616 7559 31633 7577
rect 31691 7547 31729 7589
rect 31741 7559 31758 7577
rect 31791 7559 31808 7577
rect 1281 7500 1298 7517
rect 1340 7500 1357 7517
rect 1595 7500 1612 7517
rect 1654 7500 1671 7517
rect 1909 7500 1926 7517
rect 1968 7500 1985 7517
rect 2223 7500 2240 7517
rect 2282 7500 2299 7517
rect 2537 7500 2554 7517
rect 2596 7500 2613 7517
rect 10336 7509 10380 7510
rect 9958 7486 9975 7503
rect 10017 7486 10034 7503
rect 10336 7487 10337 7509
rect 10379 7487 10380 7509
rect 12796 7509 12840 7510
rect 10668 7486 10685 7503
rect 10727 7486 10744 7503
rect 10786 7486 10803 7503
rect 11041 7486 11058 7503
rect 11100 7486 11117 7503
rect 12213 7486 12230 7503
rect 12272 7486 12289 7503
rect 12331 7486 12348 7503
rect 12586 7486 12603 7503
rect 12645 7486 12662 7503
rect 12796 7487 12797 7509
rect 12839 7487 12840 7509
rect 14600 7509 14644 7510
rect 12907 7486 12924 7503
rect 12966 7486 12983 7503
rect 13025 7486 13042 7503
rect 14600 7487 14601 7509
rect 14643 7487 14644 7509
rect 10836 7454 10846 7471
rect 12381 7454 12391 7471
rect 13075 7454 13085 7471
rect 10819 7453 10846 7454
rect 12364 7453 12391 7454
rect 13058 7453 13085 7454
rect 10757 7432 10758 7447
rect 12302 7432 12303 7447
rect 12996 7432 12997 7447
rect 13280 7444 13297 7461
rect 13349 7444 13366 7461
rect 13427 7444 13444 7461
rect 13505 7444 13522 7461
rect 13583 7444 13600 7461
rect 13661 7444 13678 7461
rect 13739 7444 13756 7461
rect 13817 7444 13834 7461
rect 13885 7444 13902 7461
rect 13366 7436 13374 7437
rect 13419 7436 13452 7437
rect 13497 7436 13505 7437
rect 13522 7436 13530 7437
rect 13575 7436 13608 7437
rect 13653 7436 13661 7437
rect 13678 7436 13686 7437
rect 13731 7436 13764 7437
rect 13809 7436 13817 7437
rect 13816 7420 13817 7428
rect 13366 7419 13391 7420
rect 13402 7419 13469 7420
rect 13480 7419 13505 7420
rect 13522 7419 13547 7420
rect 13558 7419 13625 7420
rect 13636 7419 13661 7420
rect 13678 7419 13703 7420
rect 13714 7419 13781 7420
rect 13792 7419 13817 7420
rect 1357 7377 1366 7378
rect 1671 7377 1680 7378
rect 1985 7377 1994 7378
rect 2299 7377 2308 7378
rect 2613 7377 2622 7378
rect 13856 7348 13857 7363
rect 1379 7322 1434 7331
rect 1579 7322 1675 7340
rect 1693 7322 1748 7331
rect 1893 7322 1989 7340
rect 2007 7322 2062 7331
rect 2207 7322 2303 7340
rect 2321 7322 2376 7331
rect 2521 7322 2617 7340
rect 2635 7322 2690 7331
rect 10018 7312 10034 7329
rect 11101 7312 11117 7329
rect 10018 7311 10051 7312
rect 11101 7311 11134 7312
rect 13591 7302 13600 7319
rect 13591 7301 13617 7302
rect 1281 7222 1298 7239
rect 1340 7222 1357 7239
rect 1595 7222 1612 7239
rect 1644 7221 1645 7243
rect 1654 7222 1671 7239
rect 1687 7221 1688 7243
rect 1909 7222 1926 7239
rect 1968 7222 1985 7239
rect 2223 7222 2240 7239
rect 2282 7222 2299 7239
rect 2537 7222 2554 7239
rect 2596 7222 2613 7239
rect 1644 7220 1688 7221
rect 10772 7196 10773 7211
rect 12317 7196 12318 7211
rect 12740 7203 12745 7219
rect 12723 7186 12728 7202
rect 13011 7196 13012 7211
rect 13871 7196 13872 7211
rect 1146 7185 1273 7186
rect 1306 7185 1390 7186
rect 1423 7185 1587 7186
rect 1620 7185 1704 7186
rect 1737 7185 1901 7186
rect 1934 7185 2018 7186
rect 2051 7185 2215 7186
rect 2248 7185 2332 7186
rect 2365 7185 2529 7186
rect 2562 7185 2646 7186
rect 2679 7185 2716 7186
rect 2464 7181 2508 7182
rect 2464 7159 2465 7181
rect 2507 7159 2508 7181
rect 13833 7175 13834 7183
rect 13402 7166 13468 7167
rect 13558 7166 13624 7167
rect 13714 7166 13780 7167
rect 13419 7149 13451 7150
rect 13575 7149 13607 7150
rect 13731 7149 13763 7150
rect 1281 7115 1298 7132
rect 1340 7115 1357 7132
rect 1595 7115 1612 7132
rect 1654 7115 1671 7132
rect 1909 7115 1926 7132
rect 1968 7115 1985 7132
rect 2223 7115 2240 7132
rect 2282 7115 2299 7132
rect 2537 7115 2554 7132
rect 2596 7115 2613 7132
rect 10668 7124 10685 7141
rect 10786 7124 10803 7141
rect 12213 7124 12230 7141
rect 12331 7124 12348 7141
rect 12907 7124 12924 7141
rect 13025 7124 13042 7141
rect 13280 7124 13297 7141
rect 13349 7124 13366 7141
rect 13427 7124 13444 7141
rect 13505 7124 13522 7141
rect 13583 7124 13600 7141
rect 13661 7124 13678 7141
rect 13739 7124 13756 7141
rect 13817 7124 13834 7141
rect 13885 7124 13902 7141
rect 9958 7104 9975 7121
rect 10017 7104 10034 7121
rect 11041 7104 11058 7121
rect 11100 7104 11117 7121
rect 12586 7104 12603 7121
rect 12645 7104 12662 7121
rect 12078 7067 12205 7068
rect 12238 7067 12381 7068
rect 12414 7067 12578 7068
rect 12611 7067 12695 7068
rect 12728 7067 12764 7068
rect 12781 7067 12899 7068
rect 12932 7067 13075 7068
rect 13108 7067 13272 7068
rect 13305 7067 13419 7068
rect 13451 7067 13575 7068
rect 13607 7067 13731 7068
rect 13763 7067 13877 7068
rect 13910 7067 13935 7068
rect 13944 7057 13945 7079
rect 13987 7068 13988 7079
rect 14531 7068 14569 7079
rect 31691 7068 31729 7079
rect 13968 7067 13997 7068
rect 13987 7057 13988 7067
rect 13944 7056 13988 7057
rect 14441 7050 14458 7068
rect 14534 7050 14551 7068
rect 14605 7050 14622 7068
rect 14701 7050 14718 7068
rect 14794 7050 14811 7068
rect 14865 7050 14882 7068
rect 14961 7050 14978 7068
rect 15054 7050 15071 7068
rect 15125 7050 15142 7068
rect 15221 7050 15238 7068
rect 15314 7050 15331 7068
rect 15385 7050 15402 7068
rect 15481 7050 15498 7068
rect 15574 7050 15591 7068
rect 15645 7050 15662 7068
rect 15741 7050 15758 7068
rect 15834 7050 15851 7068
rect 15905 7050 15922 7068
rect 16001 7050 16018 7068
rect 16094 7050 16111 7068
rect 16165 7050 16182 7068
rect 16261 7050 16278 7068
rect 16354 7050 16371 7068
rect 16425 7050 16442 7068
rect 16521 7050 16538 7068
rect 16614 7050 16631 7068
rect 16685 7050 16702 7068
rect 16781 7050 16798 7068
rect 16874 7050 16891 7068
rect 16945 7050 16962 7068
rect 17041 7050 17058 7068
rect 17134 7050 17151 7068
rect 17205 7050 17222 7068
rect 17301 7050 17318 7068
rect 17394 7050 17411 7068
rect 17465 7050 17482 7068
rect 17561 7050 17578 7068
rect 17654 7050 17671 7068
rect 17725 7050 17742 7068
rect 17821 7050 17838 7068
rect 17914 7050 17931 7068
rect 17985 7050 18002 7068
rect 18081 7050 18098 7068
rect 18174 7050 18191 7068
rect 18245 7050 18262 7068
rect 18341 7050 18358 7068
rect 18434 7050 18451 7068
rect 18505 7050 18522 7068
rect 18601 7050 18618 7068
rect 18694 7050 18711 7068
rect 18765 7050 18782 7068
rect 18861 7050 18878 7068
rect 18954 7050 18971 7068
rect 19025 7050 19042 7068
rect 19121 7050 19138 7068
rect 19214 7050 19231 7068
rect 19285 7050 19302 7068
rect 19381 7050 19398 7068
rect 19474 7050 19491 7068
rect 19545 7050 19562 7068
rect 19641 7050 19658 7068
rect 19734 7050 19751 7068
rect 19805 7050 19822 7068
rect 19901 7050 19918 7068
rect 19994 7050 20011 7068
rect 20065 7050 20082 7068
rect 20161 7050 20178 7068
rect 20254 7050 20271 7068
rect 20325 7050 20342 7068
rect 20421 7050 20438 7068
rect 20514 7050 20531 7068
rect 20585 7050 20602 7068
rect 20681 7050 20698 7068
rect 20774 7050 20791 7068
rect 20845 7050 20862 7068
rect 20941 7050 20958 7068
rect 21034 7050 21051 7068
rect 21105 7050 21122 7068
rect 21201 7050 21218 7068
rect 21294 7050 21311 7068
rect 21365 7050 21382 7068
rect 21461 7050 21478 7068
rect 21554 7050 21571 7068
rect 21625 7050 21642 7068
rect 21721 7050 21738 7068
rect 21814 7050 21831 7068
rect 21885 7050 21902 7068
rect 21981 7050 21998 7068
rect 22074 7050 22091 7068
rect 22145 7050 22162 7068
rect 22241 7050 22258 7068
rect 22334 7050 22351 7068
rect 22405 7050 22422 7068
rect 22501 7050 22518 7068
rect 22594 7050 22611 7068
rect 22665 7050 22682 7068
rect 22761 7050 22778 7068
rect 22854 7050 22871 7068
rect 22925 7050 22942 7068
rect 23021 7050 23038 7068
rect 23114 7050 23131 7068
rect 23185 7050 23202 7068
rect 23281 7050 23298 7068
rect 23374 7050 23391 7068
rect 23445 7050 23462 7068
rect 23541 7050 23558 7068
rect 23634 7050 23651 7068
rect 23705 7050 23722 7068
rect 23801 7050 23818 7068
rect 23894 7050 23911 7068
rect 23965 7050 23982 7068
rect 24061 7050 24078 7068
rect 24154 7050 24171 7068
rect 24225 7050 24242 7068
rect 24321 7050 24338 7068
rect 24414 7050 24431 7068
rect 24485 7050 24502 7068
rect 24581 7050 24598 7068
rect 24674 7050 24691 7068
rect 24745 7050 24762 7068
rect 24841 7050 24858 7068
rect 24934 7050 24951 7068
rect 25005 7050 25022 7068
rect 25101 7050 25118 7068
rect 25194 7050 25211 7068
rect 25265 7050 25282 7068
rect 25361 7050 25378 7068
rect 25454 7050 25471 7068
rect 25525 7050 25542 7068
rect 25621 7050 25638 7068
rect 25714 7050 25731 7068
rect 25785 7050 25802 7068
rect 25881 7050 25898 7068
rect 25974 7050 25991 7068
rect 26045 7050 26062 7068
rect 26141 7050 26158 7068
rect 26234 7050 26251 7068
rect 26305 7050 26322 7068
rect 26401 7050 26418 7068
rect 26494 7050 26511 7068
rect 26565 7050 26582 7068
rect 26661 7050 26678 7068
rect 26754 7050 26771 7068
rect 26825 7050 26842 7068
rect 26921 7050 26938 7068
rect 27014 7050 27031 7068
rect 27085 7050 27102 7068
rect 27181 7050 27198 7068
rect 27274 7050 27291 7068
rect 27345 7050 27362 7068
rect 27441 7050 27458 7068
rect 27534 7050 27551 7068
rect 27605 7050 27622 7068
rect 27701 7050 27718 7068
rect 27794 7050 27811 7068
rect 27865 7050 27882 7068
rect 27961 7050 27978 7068
rect 28054 7050 28071 7068
rect 28125 7050 28142 7068
rect 28221 7050 28238 7068
rect 28314 7050 28331 7068
rect 28385 7050 28402 7068
rect 28481 7050 28498 7068
rect 28574 7050 28591 7068
rect 28645 7050 28662 7068
rect 28741 7050 28758 7068
rect 28834 7050 28851 7068
rect 28905 7050 28922 7068
rect 29001 7050 29018 7068
rect 29094 7050 29111 7068
rect 29165 7050 29182 7068
rect 29261 7050 29278 7068
rect 29354 7050 29371 7068
rect 29425 7050 29442 7068
rect 29521 7050 29538 7068
rect 29614 7050 29631 7068
rect 29685 7050 29702 7068
rect 29781 7050 29798 7068
rect 29874 7050 29891 7068
rect 29945 7050 29962 7068
rect 30041 7050 30058 7068
rect 30134 7050 30151 7068
rect 30205 7050 30222 7068
rect 30301 7050 30318 7068
rect 30394 7050 30411 7068
rect 30465 7050 30482 7068
rect 30561 7050 30578 7068
rect 30654 7050 30671 7068
rect 30725 7050 30742 7068
rect 30821 7050 30838 7068
rect 30914 7050 30931 7068
rect 30985 7050 31002 7068
rect 31081 7050 31098 7068
rect 31174 7050 31191 7068
rect 31245 7050 31262 7068
rect 31341 7050 31358 7068
rect 31434 7050 31451 7068
rect 31505 7050 31522 7068
rect 31601 7050 31618 7068
rect 31694 7050 31711 7068
rect 31765 7050 31782 7068
rect 14531 7039 14569 7050
rect 31691 7039 31729 7050
rect 1379 7023 1434 7032
rect 1579 7014 1675 7032
rect 1693 7023 1748 7032
rect 1893 7014 1989 7032
rect 2007 7023 2062 7032
rect 2207 7014 2303 7032
rect 2321 7023 2376 7032
rect 2521 7014 2617 7032
rect 2635 7023 2690 7032
rect 10254 7017 10298 7018
rect 10254 6995 10255 7017
rect 10297 6995 10298 7017
rect 14272 7017 14316 7018
rect 14272 6995 14273 7017
rect 14315 6995 14316 7017
rect 1357 6993 1366 6994
rect 1671 6993 1680 6994
rect 1985 6993 1994 6994
rect 2299 6993 2308 6994
rect 2613 6993 2622 6994
rect 12907 6977 12924 6994
rect 13025 6977 13042 6994
rect 13280 6977 13297 6994
rect 13349 6977 13366 6994
rect 13427 6977 13444 6994
rect 13505 6977 13522 6994
rect 13583 6977 13600 6994
rect 13661 6977 13678 6994
rect 13739 6977 13756 6994
rect 13817 6977 13834 6994
rect 13885 6977 13902 6994
rect 13419 6968 13451 6969
rect 13575 6968 13607 6969
rect 13731 6968 13763 6969
rect 13816 6952 13817 6960
rect 13402 6951 13468 6952
rect 13558 6951 13624 6952
rect 13714 6951 13780 6952
rect 12996 6922 12997 6937
rect 13856 6922 13857 6937
rect 1281 6837 1298 6854
rect 1340 6837 1357 6854
rect 1595 6837 1612 6854
rect 1654 6837 1671 6854
rect 1909 6837 1926 6854
rect 1968 6837 1985 6854
rect 2223 6837 2240 6854
rect 2282 6837 2299 6854
rect 2537 6837 2554 6854
rect 2596 6837 2613 6854
rect 13591 6834 13600 6851
rect 13591 6833 13617 6834
rect 2300 6811 2301 6833
rect 2343 6811 2344 6833
rect 2300 6810 2344 6811
rect 1146 6779 1273 6780
rect 1306 6779 1390 6780
rect 1423 6779 1587 6780
rect 1620 6779 1704 6780
rect 1737 6779 1901 6780
rect 1934 6779 2018 6780
rect 2051 6779 2215 6780
rect 2248 6779 2332 6780
rect 2365 6779 2529 6780
rect 2562 6779 2646 6780
rect 2679 6779 2716 6780
rect 13871 6770 13872 6785
rect 13833 6707 13834 6715
rect 1281 6688 1298 6705
rect 1340 6688 1357 6705
rect 1595 6688 1612 6705
rect 1654 6688 1671 6705
rect 1909 6688 1926 6705
rect 1968 6688 1985 6705
rect 2223 6688 2240 6705
rect 2282 6688 2299 6705
rect 2537 6688 2554 6705
rect 2596 6688 2613 6705
rect 13011 6686 13012 6701
rect 13366 6698 13391 6699
rect 13402 6698 13469 6699
rect 13480 6698 13505 6699
rect 13522 6698 13547 6699
rect 13558 6698 13625 6699
rect 13636 6698 13661 6699
rect 13678 6698 13703 6699
rect 13714 6698 13781 6699
rect 13792 6698 13817 6699
rect 13051 6681 13059 6682
rect 13366 6681 13374 6682
rect 13419 6681 13452 6682
rect 13497 6681 13505 6682
rect 13522 6681 13530 6682
rect 13575 6681 13608 6682
rect 13653 6681 13661 6682
rect 13678 6681 13686 6682
rect 13731 6681 13764 6682
rect 13809 6681 13817 6682
rect 13058 6664 13068 6665
rect 13075 6647 13085 6665
rect 13280 6657 13297 6674
rect 13349 6657 13366 6674
rect 13427 6657 13444 6674
rect 13505 6657 13522 6674
rect 13583 6657 13600 6674
rect 13661 6657 13678 6674
rect 13739 6657 13756 6674
rect 13817 6657 13834 6674
rect 13885 6657 13902 6674
rect 12907 6615 12924 6632
rect 12966 6615 12983 6632
rect 13025 6615 13042 6632
rect 1357 6565 1366 6566
rect 1671 6565 1680 6566
rect 1985 6565 1994 6566
rect 2299 6565 2308 6566
rect 2613 6565 2622 6566
rect 14456 6541 14473 6559
rect 14531 6529 14569 6571
rect 14581 6541 14598 6559
rect 14631 6541 14648 6559
rect 14716 6541 14733 6559
rect 14794 6541 14811 6559
rect 14841 6541 14858 6559
rect 14891 6541 14908 6559
rect 14976 6541 14993 6559
rect 15054 6541 15071 6559
rect 15101 6541 15118 6559
rect 15151 6541 15168 6559
rect 15236 6541 15253 6559
rect 15314 6541 15331 6559
rect 15361 6541 15378 6559
rect 15411 6541 15428 6559
rect 15496 6541 15513 6559
rect 15574 6541 15591 6559
rect 15621 6541 15638 6559
rect 15671 6541 15688 6559
rect 15756 6541 15773 6559
rect 15834 6541 15851 6559
rect 15881 6541 15898 6559
rect 15931 6541 15948 6559
rect 16016 6541 16033 6559
rect 16094 6541 16111 6559
rect 16141 6541 16158 6559
rect 16191 6541 16208 6559
rect 16276 6541 16293 6559
rect 16354 6541 16371 6559
rect 16401 6541 16418 6559
rect 16451 6541 16468 6559
rect 16536 6541 16553 6559
rect 16614 6541 16631 6559
rect 16661 6541 16678 6559
rect 16711 6541 16728 6559
rect 16796 6541 16813 6559
rect 16874 6541 16891 6559
rect 16921 6541 16938 6559
rect 16971 6541 16988 6559
rect 17056 6541 17073 6559
rect 17134 6541 17151 6559
rect 17181 6541 17198 6559
rect 17231 6541 17248 6559
rect 17316 6541 17333 6559
rect 17394 6541 17411 6559
rect 17441 6541 17458 6559
rect 17491 6541 17508 6559
rect 17576 6541 17593 6559
rect 17654 6541 17671 6559
rect 17701 6541 17718 6559
rect 17751 6541 17768 6559
rect 17836 6541 17853 6559
rect 17914 6541 17931 6559
rect 17961 6541 17978 6559
rect 18011 6541 18028 6559
rect 18096 6541 18113 6559
rect 18174 6541 18191 6559
rect 18221 6541 18238 6559
rect 18271 6541 18288 6559
rect 18356 6541 18373 6559
rect 18434 6541 18451 6559
rect 18481 6541 18498 6559
rect 18531 6541 18548 6559
rect 18616 6541 18633 6559
rect 18694 6541 18711 6559
rect 18741 6541 18758 6559
rect 18791 6541 18808 6559
rect 18876 6541 18893 6559
rect 18954 6541 18971 6559
rect 19001 6541 19018 6559
rect 19051 6541 19068 6559
rect 19136 6541 19153 6559
rect 19214 6541 19231 6559
rect 19261 6541 19278 6559
rect 19311 6541 19328 6559
rect 19396 6541 19413 6559
rect 19474 6541 19491 6559
rect 19521 6541 19538 6559
rect 19571 6541 19588 6559
rect 19656 6541 19673 6559
rect 19734 6541 19751 6559
rect 19781 6541 19798 6559
rect 19831 6541 19848 6559
rect 19916 6541 19933 6559
rect 19994 6541 20011 6559
rect 20041 6541 20058 6559
rect 20091 6541 20108 6559
rect 20176 6541 20193 6559
rect 20254 6541 20271 6559
rect 20301 6541 20318 6559
rect 20351 6541 20368 6559
rect 20436 6541 20453 6559
rect 20514 6541 20531 6559
rect 20561 6541 20578 6559
rect 20611 6541 20628 6559
rect 20696 6541 20713 6559
rect 20774 6541 20791 6559
rect 20821 6541 20838 6559
rect 20871 6541 20888 6559
rect 20956 6541 20973 6559
rect 21034 6541 21051 6559
rect 21081 6541 21098 6559
rect 21131 6541 21148 6559
rect 21216 6541 21233 6559
rect 21294 6541 21311 6559
rect 21341 6541 21358 6559
rect 21391 6541 21408 6559
rect 21476 6541 21493 6559
rect 21554 6541 21571 6559
rect 21601 6541 21618 6559
rect 21651 6541 21668 6559
rect 21736 6541 21753 6559
rect 21814 6541 21831 6559
rect 21861 6541 21878 6559
rect 21911 6541 21928 6559
rect 21996 6541 22013 6559
rect 22074 6541 22091 6559
rect 22121 6541 22138 6559
rect 22171 6541 22188 6559
rect 22256 6541 22273 6559
rect 22334 6541 22351 6559
rect 22381 6541 22398 6559
rect 22431 6541 22448 6559
rect 22516 6541 22533 6559
rect 22594 6541 22611 6559
rect 22641 6541 22658 6559
rect 22691 6541 22708 6559
rect 22776 6541 22793 6559
rect 22854 6541 22871 6559
rect 22901 6541 22918 6559
rect 22951 6541 22968 6559
rect 23036 6541 23053 6559
rect 23114 6541 23131 6559
rect 23161 6541 23178 6559
rect 23211 6541 23228 6559
rect 23296 6541 23313 6559
rect 23374 6541 23391 6559
rect 23421 6541 23438 6559
rect 23471 6541 23488 6559
rect 23556 6541 23573 6559
rect 23634 6541 23651 6559
rect 23681 6541 23698 6559
rect 23731 6541 23748 6559
rect 23816 6541 23833 6559
rect 23894 6541 23911 6559
rect 23941 6541 23958 6559
rect 23991 6541 24008 6559
rect 24076 6541 24093 6559
rect 24154 6541 24171 6559
rect 24201 6541 24218 6559
rect 24251 6541 24268 6559
rect 24336 6541 24353 6559
rect 24414 6541 24431 6559
rect 24461 6541 24478 6559
rect 24511 6541 24528 6559
rect 24596 6541 24613 6559
rect 24674 6541 24691 6559
rect 24721 6541 24738 6559
rect 24771 6541 24788 6559
rect 24856 6541 24873 6559
rect 24934 6541 24951 6559
rect 24981 6541 24998 6559
rect 25031 6541 25048 6559
rect 25116 6541 25133 6559
rect 25194 6541 25211 6559
rect 25241 6541 25258 6559
rect 25291 6541 25308 6559
rect 25376 6541 25393 6559
rect 25454 6541 25471 6559
rect 25501 6541 25518 6559
rect 25551 6541 25568 6559
rect 25636 6541 25653 6559
rect 25714 6541 25731 6559
rect 25761 6541 25778 6559
rect 25811 6541 25828 6559
rect 25896 6541 25913 6559
rect 25974 6541 25991 6559
rect 26021 6541 26038 6559
rect 26071 6541 26088 6559
rect 26156 6541 26173 6559
rect 26234 6541 26251 6559
rect 26281 6541 26298 6559
rect 26331 6541 26348 6559
rect 26416 6541 26433 6559
rect 26494 6541 26511 6559
rect 26541 6541 26558 6559
rect 26591 6541 26608 6559
rect 26676 6541 26693 6559
rect 26754 6541 26771 6559
rect 26801 6541 26818 6559
rect 26851 6541 26868 6559
rect 26936 6541 26953 6559
rect 27014 6541 27031 6559
rect 27061 6541 27078 6559
rect 27111 6541 27128 6559
rect 27196 6541 27213 6559
rect 27274 6541 27291 6559
rect 27321 6541 27338 6559
rect 27371 6541 27388 6559
rect 27456 6541 27473 6559
rect 27534 6541 27551 6559
rect 27581 6541 27598 6559
rect 27631 6541 27648 6559
rect 27716 6541 27733 6559
rect 27794 6541 27811 6559
rect 27841 6541 27858 6559
rect 27891 6541 27908 6559
rect 27976 6541 27993 6559
rect 28054 6541 28071 6559
rect 28101 6541 28118 6559
rect 28151 6541 28168 6559
rect 28236 6541 28253 6559
rect 28314 6541 28331 6559
rect 28361 6541 28378 6559
rect 28411 6541 28428 6559
rect 28496 6541 28513 6559
rect 28574 6541 28591 6559
rect 28621 6541 28638 6559
rect 28671 6541 28688 6559
rect 28756 6541 28773 6559
rect 28834 6541 28851 6559
rect 28881 6541 28898 6559
rect 28931 6541 28948 6559
rect 29016 6541 29033 6559
rect 29094 6541 29111 6559
rect 29141 6541 29158 6559
rect 29191 6541 29208 6559
rect 29276 6541 29293 6559
rect 29354 6541 29371 6559
rect 29401 6541 29418 6559
rect 29451 6541 29468 6559
rect 29536 6541 29553 6559
rect 29614 6541 29631 6559
rect 29661 6541 29678 6559
rect 29711 6541 29728 6559
rect 29796 6541 29813 6559
rect 29874 6541 29891 6559
rect 29921 6541 29938 6559
rect 29971 6541 29988 6559
rect 30056 6541 30073 6559
rect 30134 6541 30151 6559
rect 30181 6541 30198 6559
rect 30231 6541 30248 6559
rect 30316 6541 30333 6559
rect 30394 6541 30411 6559
rect 30441 6541 30458 6559
rect 30491 6541 30508 6559
rect 30576 6541 30593 6559
rect 30654 6541 30671 6559
rect 30701 6541 30718 6559
rect 30751 6541 30768 6559
rect 30836 6541 30853 6559
rect 30914 6541 30931 6559
rect 30961 6541 30978 6559
rect 31011 6541 31028 6559
rect 31096 6541 31113 6559
rect 31174 6541 31191 6559
rect 31221 6541 31238 6559
rect 31271 6541 31288 6559
rect 31356 6541 31373 6559
rect 31434 6541 31451 6559
rect 31481 6541 31498 6559
rect 31531 6541 31548 6559
rect 31616 6541 31633 6559
rect 31691 6529 31729 6571
rect 31741 6541 31758 6559
rect 31791 6541 31808 6559
rect 1379 6510 1434 6519
rect 1579 6510 1675 6528
rect 1693 6510 1748 6519
rect 1893 6510 1989 6528
rect 2007 6510 2062 6519
rect 2207 6510 2303 6528
rect 2321 6510 2376 6519
rect 2521 6510 2617 6528
rect 14682 6525 14726 6526
rect 2635 6510 2690 6519
rect 14682 6503 14683 6525
rect 14725 6503 14726 6525
rect 1281 6410 1298 6427
rect 1340 6410 1357 6427
rect 1595 6410 1612 6427
rect 1654 6410 1671 6427
rect 1909 6410 1926 6427
rect 1968 6410 1985 6427
rect 2223 6410 2240 6427
rect 2282 6410 2299 6427
rect 2537 6410 2554 6427
rect 2596 6410 2613 6427
rect 1146 6373 1273 6374
rect 1306 6373 1390 6374
rect 1423 6373 1587 6374
rect 1620 6373 1704 6374
rect 1737 6373 1901 6374
rect 1934 6373 2018 6374
rect 2051 6373 2215 6374
rect 2248 6373 2332 6374
rect 2365 6373 2529 6374
rect 2562 6373 2646 6374
rect 2679 6373 2716 6374
rect 1281 6303 1298 6320
rect 1340 6303 1357 6320
rect 1595 6303 1612 6320
rect 1654 6303 1671 6320
rect 1909 6303 1926 6320
rect 1968 6303 1985 6320
rect 2223 6303 2240 6320
rect 2282 6303 2299 6320
rect 2537 6303 2554 6320
rect 2596 6303 2613 6320
rect 1379 6211 1434 6220
rect 1579 6202 1675 6220
rect 1693 6211 1748 6220
rect 1893 6202 1989 6220
rect 2007 6211 2062 6220
rect 2207 6202 2303 6220
rect 2321 6211 2376 6220
rect 2521 6202 2617 6220
rect 2635 6211 2690 6220
rect 1357 6181 1366 6182
rect 1671 6181 1680 6182
rect 1985 6181 1994 6182
rect 2299 6181 2308 6182
rect 2613 6181 2622 6182
rect 31492 6073 31493 6095
rect 31535 6073 31536 6095
rect 31492 6072 31536 6073
rect 1281 6025 1298 6042
rect 1340 6025 1357 6042
rect 1595 6025 1612 6042
rect 1654 6025 1671 6042
rect 1909 6025 1926 6042
rect 1968 6025 1985 6042
rect 2223 6025 2240 6042
rect 2282 6025 2299 6042
rect 2537 6025 2554 6042
rect 2596 6025 2613 6042
rect 14745 6021 14747 6041
rect 2382 5991 2383 6013
rect 2425 5991 2426 6013
rect 14759 6007 14761 6041
rect 14770 6001 14773 6041
rect 14784 6015 14787 6041
rect 14832 6015 14836 6041
rect 14846 6001 14850 6041
rect 15005 6021 15007 6041
rect 15019 6007 15021 6041
rect 15030 6001 15033 6041
rect 15044 6015 15047 6041
rect 15092 6015 15096 6041
rect 15106 6001 15110 6041
rect 15265 6021 15267 6041
rect 15279 6007 15281 6041
rect 15290 6001 15293 6041
rect 15304 6015 15307 6041
rect 15352 6015 15356 6041
rect 15366 6001 15370 6041
rect 15525 6021 15527 6041
rect 15539 6007 15541 6041
rect 15550 6001 15553 6041
rect 15564 6015 15567 6041
rect 15612 6015 15616 6041
rect 15626 6001 15630 6041
rect 15785 6021 15787 6041
rect 15799 6007 15801 6041
rect 15810 6001 15813 6041
rect 15824 6015 15827 6041
rect 15872 6015 15876 6041
rect 15886 6001 15890 6041
rect 16045 6021 16047 6041
rect 16059 6007 16061 6041
rect 16070 6001 16073 6041
rect 16084 6015 16087 6041
rect 16132 6015 16136 6041
rect 16146 6001 16150 6041
rect 16305 6021 16307 6041
rect 16319 6007 16321 6041
rect 16330 6001 16333 6041
rect 16344 6015 16347 6041
rect 16392 6015 16396 6041
rect 16406 6001 16410 6041
rect 16565 6021 16567 6041
rect 16579 6007 16581 6041
rect 16590 6001 16593 6041
rect 16604 6015 16607 6041
rect 16652 6015 16656 6041
rect 16666 6001 16670 6041
rect 16825 6021 16827 6041
rect 16839 6007 16841 6041
rect 16850 6001 16853 6041
rect 16864 6015 16867 6041
rect 16912 6015 16916 6041
rect 16926 6001 16930 6041
rect 17085 6021 17087 6041
rect 17099 6007 17101 6041
rect 17110 6001 17113 6041
rect 17124 6015 17127 6041
rect 17172 6015 17176 6041
rect 17186 6001 17190 6041
rect 17345 6021 17347 6041
rect 17359 6007 17361 6041
rect 17370 6001 17373 6041
rect 17384 6015 17387 6041
rect 17432 6015 17436 6041
rect 17446 6001 17450 6041
rect 17605 6021 17607 6041
rect 17619 6007 17621 6041
rect 17630 6001 17633 6041
rect 17644 6015 17647 6041
rect 17692 6015 17696 6041
rect 17706 6001 17710 6041
rect 17865 6021 17867 6041
rect 17879 6007 17881 6041
rect 17890 6001 17893 6041
rect 17904 6015 17907 6041
rect 17952 6015 17956 6041
rect 17966 6001 17970 6041
rect 18125 6021 18127 6041
rect 18139 6007 18141 6041
rect 18150 6001 18153 6041
rect 18164 6015 18167 6041
rect 18212 6015 18216 6041
rect 18226 6001 18230 6041
rect 18385 6021 18387 6041
rect 18399 6007 18401 6041
rect 18410 6001 18413 6041
rect 18424 6015 18427 6041
rect 18472 6015 18476 6041
rect 18486 6001 18490 6041
rect 18645 6021 18647 6041
rect 18659 6007 18661 6041
rect 18670 6001 18673 6041
rect 18684 6015 18687 6041
rect 18732 6015 18736 6041
rect 18746 6001 18750 6041
rect 18905 6021 18907 6041
rect 18919 6007 18921 6041
rect 18930 6001 18933 6041
rect 18944 6015 18947 6041
rect 18992 6015 18996 6041
rect 19006 6001 19010 6041
rect 19165 6021 19167 6041
rect 19179 6007 19181 6041
rect 19190 6001 19193 6041
rect 19204 6015 19207 6041
rect 19252 6015 19256 6041
rect 19266 6001 19270 6041
rect 19425 6021 19427 6041
rect 19439 6007 19441 6041
rect 19450 6001 19453 6041
rect 19464 6015 19467 6041
rect 19512 6015 19516 6041
rect 19526 6001 19530 6041
rect 19685 6021 19687 6041
rect 19699 6007 19701 6041
rect 19710 6001 19713 6041
rect 19724 6015 19727 6041
rect 19772 6015 19776 6041
rect 19786 6001 19790 6041
rect 19945 6021 19947 6041
rect 19959 6007 19961 6041
rect 19970 6001 19973 6041
rect 19984 6015 19987 6041
rect 20032 6015 20036 6041
rect 20046 6001 20050 6041
rect 20205 6021 20207 6041
rect 20219 6007 20221 6041
rect 20230 6001 20233 6041
rect 20244 6015 20247 6041
rect 20292 6015 20296 6041
rect 20306 6001 20310 6041
rect 20465 6021 20467 6041
rect 20479 6007 20481 6041
rect 20490 6001 20493 6041
rect 20504 6015 20507 6041
rect 20552 6015 20556 6041
rect 20566 6001 20570 6041
rect 20725 6021 20727 6041
rect 20739 6007 20741 6041
rect 20750 6001 20753 6041
rect 20764 6015 20767 6041
rect 20812 6015 20816 6041
rect 20826 6001 20830 6041
rect 20985 6021 20987 6041
rect 20999 6007 21001 6041
rect 21010 6001 21013 6041
rect 21024 6015 21027 6041
rect 21072 6015 21076 6041
rect 21086 6001 21090 6041
rect 21245 6021 21247 6041
rect 21259 6007 21261 6041
rect 21270 6001 21273 6041
rect 21284 6015 21287 6041
rect 21332 6015 21336 6041
rect 21346 6001 21350 6041
rect 21505 6021 21507 6041
rect 21519 6007 21521 6041
rect 21530 6001 21533 6041
rect 21544 6015 21547 6041
rect 21592 6015 21596 6041
rect 21606 6001 21610 6041
rect 21765 6021 21767 6041
rect 21779 6007 21781 6041
rect 21790 6001 21793 6041
rect 21804 6015 21807 6041
rect 21852 6015 21856 6041
rect 21866 6001 21870 6041
rect 22025 6021 22027 6041
rect 22039 6007 22041 6041
rect 22050 6001 22053 6041
rect 22064 6015 22067 6041
rect 22112 6015 22116 6041
rect 22126 6001 22130 6041
rect 22285 6021 22287 6041
rect 22299 6007 22301 6041
rect 22310 6001 22313 6041
rect 22324 6015 22327 6041
rect 22372 6015 22376 6041
rect 22386 6001 22390 6041
rect 22545 6021 22547 6041
rect 22559 6007 22561 6041
rect 22570 6001 22573 6041
rect 22584 6015 22587 6041
rect 22632 6015 22636 6041
rect 22646 6001 22650 6041
rect 22805 6021 22807 6041
rect 22819 6007 22821 6041
rect 22830 6001 22833 6041
rect 22844 6015 22847 6041
rect 22892 6015 22896 6041
rect 22906 6001 22910 6041
rect 23065 6021 23067 6041
rect 23079 6007 23081 6041
rect 23090 6001 23093 6041
rect 23104 6015 23107 6041
rect 23152 6015 23156 6041
rect 23166 6001 23170 6041
rect 23325 6021 23327 6041
rect 23339 6007 23341 6041
rect 23350 6001 23353 6041
rect 23364 6015 23367 6041
rect 23412 6015 23416 6041
rect 23426 6001 23430 6041
rect 23585 6021 23587 6041
rect 23599 6007 23601 6041
rect 23610 6001 23613 6041
rect 23624 6015 23627 6041
rect 23672 6015 23676 6041
rect 23686 6001 23690 6041
rect 23845 6021 23847 6041
rect 23859 6007 23861 6041
rect 23870 6001 23873 6041
rect 23884 6015 23887 6041
rect 23932 6015 23936 6041
rect 23946 6001 23950 6041
rect 24105 6021 24107 6041
rect 24119 6007 24121 6041
rect 24130 6001 24133 6041
rect 24144 6015 24147 6041
rect 24192 6015 24196 6041
rect 24206 6001 24210 6041
rect 24365 6021 24367 6041
rect 24379 6007 24381 6041
rect 24390 6001 24393 6041
rect 24404 6015 24407 6041
rect 24452 6015 24456 6041
rect 24466 6001 24470 6041
rect 24625 6021 24627 6041
rect 24639 6007 24641 6041
rect 24650 6001 24653 6041
rect 24664 6015 24667 6041
rect 24712 6015 24716 6041
rect 24726 6001 24730 6041
rect 24885 6021 24887 6041
rect 24899 6007 24901 6041
rect 24910 6001 24913 6041
rect 24924 6015 24927 6041
rect 24972 6015 24976 6041
rect 24986 6001 24990 6041
rect 25145 6021 25147 6041
rect 25159 6007 25161 6041
rect 25170 6001 25173 6041
rect 25184 6015 25187 6041
rect 25232 6015 25236 6041
rect 25246 6001 25250 6041
rect 25405 6021 25407 6041
rect 25419 6007 25421 6041
rect 25430 6001 25433 6041
rect 25444 6015 25447 6041
rect 25492 6015 25496 6041
rect 25506 6001 25510 6041
rect 25665 6021 25667 6041
rect 25679 6007 25681 6041
rect 25690 6001 25693 6041
rect 25704 6015 25707 6041
rect 25752 6015 25756 6041
rect 25766 6001 25770 6041
rect 25925 6021 25927 6041
rect 25939 6007 25941 6041
rect 25950 6001 25953 6041
rect 25964 6015 25967 6041
rect 26012 6015 26016 6041
rect 26026 6001 26030 6041
rect 26185 6021 26187 6041
rect 26199 6007 26201 6041
rect 26210 6001 26213 6041
rect 26224 6015 26227 6041
rect 26272 6015 26276 6041
rect 26286 6001 26290 6041
rect 26445 6021 26447 6041
rect 26459 6007 26461 6041
rect 26470 6001 26473 6041
rect 26484 6015 26487 6041
rect 26532 6015 26536 6041
rect 26546 6001 26550 6041
rect 26705 6021 26707 6041
rect 26719 6007 26721 6041
rect 26730 6001 26733 6041
rect 26744 6015 26747 6041
rect 26792 6015 26796 6041
rect 26806 6001 26810 6041
rect 26965 6021 26967 6041
rect 26979 6007 26981 6041
rect 26990 6001 26993 6041
rect 27004 6015 27007 6041
rect 27052 6015 27056 6041
rect 27066 6001 27070 6041
rect 27225 6021 27227 6041
rect 27239 6007 27241 6041
rect 27250 6001 27253 6041
rect 27264 6015 27267 6041
rect 27312 6015 27316 6041
rect 27326 6001 27330 6041
rect 27485 6021 27487 6041
rect 27499 6007 27501 6041
rect 27510 6001 27513 6041
rect 27524 6015 27527 6041
rect 27572 6015 27576 6041
rect 27586 6001 27590 6041
rect 27745 6021 27747 6041
rect 27759 6007 27761 6041
rect 27770 6001 27773 6041
rect 27784 6015 27787 6041
rect 27832 6015 27836 6041
rect 27846 6001 27850 6041
rect 28005 6021 28007 6041
rect 28019 6007 28021 6041
rect 28030 6001 28033 6041
rect 28044 6015 28047 6041
rect 28092 6015 28096 6041
rect 28106 6001 28110 6041
rect 28265 6021 28267 6041
rect 28279 6007 28281 6041
rect 28290 6001 28293 6041
rect 28304 6015 28307 6041
rect 28352 6015 28356 6041
rect 28366 6001 28370 6041
rect 28525 6021 28527 6041
rect 28539 6007 28541 6041
rect 28550 6001 28553 6041
rect 28564 6015 28567 6041
rect 28612 6015 28616 6041
rect 28626 6001 28630 6041
rect 28785 6021 28787 6041
rect 28799 6007 28801 6041
rect 28810 6001 28813 6041
rect 28824 6015 28827 6041
rect 28872 6015 28876 6041
rect 28886 6001 28890 6041
rect 29045 6021 29047 6041
rect 29059 6007 29061 6041
rect 29070 6001 29073 6041
rect 29084 6015 29087 6041
rect 29132 6015 29136 6041
rect 29146 6001 29150 6041
rect 29305 6021 29307 6041
rect 29319 6007 29321 6041
rect 29330 6001 29333 6041
rect 29344 6015 29347 6041
rect 29392 6015 29396 6041
rect 29406 6001 29410 6041
rect 29565 6021 29567 6041
rect 29579 6007 29581 6041
rect 29590 6001 29593 6041
rect 29604 6015 29607 6041
rect 29652 6015 29656 6041
rect 29666 6001 29670 6041
rect 29825 6021 29827 6041
rect 29839 6007 29841 6041
rect 29850 6001 29853 6041
rect 29864 6015 29867 6041
rect 29912 6015 29916 6041
rect 29926 6001 29930 6041
rect 30085 6021 30087 6041
rect 30099 6007 30101 6041
rect 30110 6001 30113 6041
rect 30124 6015 30127 6041
rect 30172 6015 30176 6041
rect 30186 6001 30190 6041
rect 30345 6021 30347 6041
rect 30359 6007 30361 6041
rect 30370 6001 30373 6041
rect 30384 6015 30387 6041
rect 30432 6015 30436 6041
rect 30446 6001 30450 6041
rect 30605 6021 30607 6041
rect 30619 6007 30621 6041
rect 30630 6001 30633 6041
rect 30644 6015 30647 6041
rect 30692 6015 30696 6041
rect 30706 6001 30710 6041
rect 30865 6021 30867 6041
rect 30879 6007 30881 6041
rect 30890 6001 30893 6041
rect 30904 6015 30907 6041
rect 30952 6015 30956 6041
rect 30966 6001 30970 6041
rect 31125 6021 31127 6041
rect 31139 6007 31141 6041
rect 31150 6001 31153 6041
rect 31164 6015 31167 6041
rect 31212 6015 31216 6041
rect 31226 6001 31230 6041
rect 31385 6021 31387 6041
rect 31399 6007 31401 6041
rect 31410 6001 31413 6041
rect 31424 6015 31427 6041
rect 31472 6015 31476 6041
rect 31486 6001 31490 6041
rect 2382 5990 2426 5991
rect 1146 5967 1273 5968
rect 1306 5967 1390 5968
rect 1423 5967 1587 5968
rect 1620 5967 1704 5968
rect 1737 5967 1901 5968
rect 1934 5967 2018 5968
rect 2051 5967 2215 5968
rect 2248 5967 2332 5968
rect 2365 5967 2529 5968
rect 2562 5967 2646 5968
rect 2679 5967 2716 5968
rect 4148 5967 5400 5968
rect 4283 5897 4300 5914
rect 4352 5897 4369 5914
rect 4430 5897 4447 5914
rect 4498 5897 4515 5914
rect 1281 5876 1298 5893
rect 1340 5876 1357 5893
rect 1595 5876 1612 5893
rect 1654 5876 1671 5893
rect 1909 5876 1926 5893
rect 1968 5876 1985 5893
rect 2223 5876 2240 5893
rect 2282 5876 2299 5893
rect 2537 5876 2554 5893
rect 2596 5876 2613 5893
rect 4753 5889 4770 5906
rect 4822 5889 4839 5906
rect 4900 5889 4917 5906
rect 4978 5889 4995 5906
rect 5056 5889 5073 5906
rect 5134 5889 5151 5906
rect 5212 5889 5229 5906
rect 5280 5889 5297 5906
rect 4892 5880 4924 5881
rect 5048 5880 5080 5881
rect 5204 5880 5236 5881
rect 4469 5873 4470 5879
rect 4369 5872 4498 5873
rect 4469 5864 4470 5872
rect 4875 5863 4941 5864
rect 5031 5863 5097 5864
rect 5187 5863 5253 5864
rect 5251 5846 5252 5861
rect 4537 5805 4592 5814
rect 5319 5805 5374 5832
rect 1357 5753 1366 5754
rect 1671 5753 1680 5754
rect 1985 5753 1994 5754
rect 2299 5753 2308 5754
rect 2613 5753 2622 5754
rect 5266 5726 5267 5741
rect 1379 5698 1434 5707
rect 1579 5698 1675 5716
rect 1693 5698 1748 5707
rect 1893 5698 1989 5716
rect 2007 5698 2062 5707
rect 2207 5698 2303 5716
rect 2321 5698 2376 5707
rect 2521 5698 2617 5716
rect 2635 5698 2690 5707
rect 4484 5690 4485 5705
rect 4839 5678 4864 5679
rect 4875 5678 4942 5679
rect 4953 5678 4978 5679
rect 4995 5678 5020 5679
rect 5031 5678 5098 5679
rect 5109 5678 5134 5679
rect 5151 5678 5176 5679
rect 5187 5678 5254 5679
rect 5255 5678 5280 5679
rect 4839 5661 4847 5662
rect 4892 5661 4925 5662
rect 4970 5661 4978 5662
rect 4995 5661 5003 5662
rect 5048 5661 5081 5662
rect 5126 5661 5134 5662
rect 5151 5661 5159 5662
rect 5204 5661 5237 5662
rect 5272 5661 5280 5662
rect 4369 5660 4394 5661
rect 4405 5660 4472 5661
rect 4473 5660 4498 5661
rect 4369 5643 4377 5644
rect 4422 5643 4455 5644
rect 4490 5643 4498 5644
rect 4753 5637 4770 5654
rect 4822 5637 4839 5654
rect 4900 5637 4917 5654
rect 4978 5637 4995 5654
rect 5056 5637 5073 5654
rect 5134 5637 5151 5654
rect 5212 5637 5229 5654
rect 5280 5637 5297 5654
rect 4283 5619 4300 5636
rect 4352 5619 4369 5636
rect 4430 5619 4447 5636
rect 4498 5619 4515 5636
rect 1281 5598 1298 5615
rect 1340 5598 1357 5615
rect 1595 5598 1612 5615
rect 1654 5598 1671 5615
rect 1726 5581 1727 5603
rect 1769 5581 1770 5603
rect 1909 5598 1926 5615
rect 1968 5598 1985 5615
rect 2223 5598 2240 5615
rect 2282 5598 2299 5615
rect 2537 5598 2554 5615
rect 2596 5598 2613 5615
rect 14822 5585 14839 5602
rect 1726 5580 1770 5581
rect 14853 5571 14854 5617
rect 1146 5561 1273 5562
rect 1306 5561 1390 5562
rect 1423 5561 1587 5562
rect 1620 5561 1704 5562
rect 1737 5561 1901 5562
rect 1934 5561 2018 5562
rect 2051 5561 2215 5562
rect 2248 5561 2332 5562
rect 2365 5561 2529 5562
rect 2562 5561 2646 5562
rect 2679 5561 2716 5562
rect 4148 5561 4275 5562
rect 4308 5561 4422 5562
rect 4454 5561 4548 5562
rect 4581 5561 4745 5562
rect 4778 5561 4892 5562
rect 4924 5561 5048 5562
rect 5080 5561 5204 5562
rect 5236 5561 5330 5562
rect 5363 5561 5400 5562
rect 14867 5557 14868 5631
rect 14881 5585 14898 5602
rect 14940 5585 14957 5602
rect 15082 5585 15099 5602
rect 15113 5571 15114 5617
rect 15127 5557 15128 5631
rect 15141 5585 15158 5602
rect 15200 5585 15217 5602
rect 15342 5585 15359 5602
rect 15373 5571 15374 5617
rect 15387 5557 15388 5631
rect 15401 5585 15418 5602
rect 15460 5585 15477 5602
rect 15602 5585 15619 5602
rect 15633 5571 15634 5617
rect 15647 5557 15648 5631
rect 15661 5585 15678 5602
rect 15720 5585 15737 5602
rect 15862 5585 15879 5602
rect 15893 5571 15894 5617
rect 15907 5557 15908 5631
rect 15921 5585 15938 5602
rect 15980 5585 15997 5602
rect 16122 5585 16139 5602
rect 16153 5571 16154 5617
rect 16167 5557 16168 5631
rect 16181 5585 16198 5602
rect 16240 5585 16257 5602
rect 16382 5585 16399 5602
rect 16413 5571 16414 5617
rect 16427 5557 16428 5631
rect 16441 5585 16458 5602
rect 16500 5585 16517 5602
rect 16642 5585 16659 5602
rect 16673 5571 16674 5617
rect 16687 5557 16688 5631
rect 16701 5585 16718 5602
rect 16760 5585 16777 5602
rect 16902 5585 16919 5602
rect 16933 5571 16934 5617
rect 16947 5557 16948 5631
rect 16961 5585 16978 5602
rect 17020 5585 17037 5602
rect 17162 5585 17179 5602
rect 17193 5571 17194 5617
rect 17207 5557 17208 5631
rect 17221 5585 17238 5602
rect 17280 5585 17297 5602
rect 17422 5585 17439 5602
rect 17453 5571 17454 5617
rect 17467 5557 17468 5631
rect 17481 5585 17498 5602
rect 17540 5585 17557 5602
rect 17682 5585 17699 5602
rect 17713 5571 17714 5617
rect 17727 5557 17728 5631
rect 17741 5585 17758 5602
rect 17800 5585 17817 5602
rect 17942 5585 17959 5602
rect 17973 5571 17974 5617
rect 17987 5557 17988 5631
rect 18001 5585 18018 5602
rect 18060 5585 18077 5602
rect 18202 5585 18219 5602
rect 18233 5571 18234 5617
rect 18247 5557 18248 5631
rect 18261 5585 18278 5602
rect 18320 5585 18337 5602
rect 18462 5585 18479 5602
rect 18493 5571 18494 5617
rect 18507 5557 18508 5631
rect 18521 5585 18538 5602
rect 18580 5585 18597 5602
rect 18722 5585 18739 5602
rect 18753 5571 18754 5617
rect 18767 5557 18768 5631
rect 18781 5585 18798 5602
rect 18840 5585 18857 5602
rect 18982 5585 18999 5602
rect 19013 5571 19014 5617
rect 19027 5557 19028 5631
rect 19041 5585 19058 5602
rect 19100 5585 19117 5602
rect 19242 5585 19259 5602
rect 19273 5571 19274 5617
rect 19287 5557 19288 5631
rect 19301 5585 19318 5602
rect 19360 5585 19377 5602
rect 19502 5585 19519 5602
rect 19533 5571 19534 5617
rect 19547 5557 19548 5631
rect 19561 5585 19578 5602
rect 19620 5585 19637 5602
rect 19762 5585 19779 5602
rect 19793 5571 19794 5617
rect 19807 5557 19808 5631
rect 19821 5585 19838 5602
rect 19880 5585 19897 5602
rect 20022 5585 20039 5602
rect 20053 5571 20054 5617
rect 20067 5557 20068 5631
rect 20081 5585 20098 5602
rect 20140 5585 20157 5602
rect 20282 5585 20299 5602
rect 20313 5571 20314 5617
rect 20327 5557 20328 5631
rect 20341 5585 20358 5602
rect 20400 5585 20417 5602
rect 20542 5585 20559 5602
rect 20573 5571 20574 5617
rect 20587 5557 20588 5631
rect 20601 5585 20618 5602
rect 20660 5585 20677 5602
rect 20802 5585 20819 5602
rect 20833 5571 20834 5617
rect 20847 5557 20848 5631
rect 20861 5585 20878 5602
rect 20920 5585 20937 5602
rect 21062 5585 21079 5602
rect 21093 5571 21094 5617
rect 21107 5557 21108 5631
rect 21121 5585 21138 5602
rect 21180 5585 21197 5602
rect 21322 5585 21339 5602
rect 21353 5571 21354 5617
rect 21367 5557 21368 5631
rect 21381 5585 21398 5602
rect 21440 5585 21457 5602
rect 21582 5585 21599 5602
rect 21613 5571 21614 5617
rect 21627 5557 21628 5631
rect 21641 5585 21658 5602
rect 21700 5585 21717 5602
rect 21842 5585 21859 5602
rect 21873 5571 21874 5617
rect 21887 5557 21888 5631
rect 21901 5585 21918 5602
rect 21960 5585 21977 5602
rect 22102 5585 22119 5602
rect 22133 5571 22134 5617
rect 22147 5557 22148 5631
rect 22161 5585 22178 5602
rect 22220 5585 22237 5602
rect 22362 5585 22379 5602
rect 22393 5571 22394 5617
rect 22407 5557 22408 5631
rect 22421 5585 22438 5602
rect 22480 5585 22497 5602
rect 22622 5585 22639 5602
rect 22653 5571 22654 5617
rect 22667 5557 22668 5631
rect 22681 5585 22698 5602
rect 22740 5585 22757 5602
rect 22882 5585 22899 5602
rect 22913 5571 22914 5617
rect 22927 5557 22928 5631
rect 22941 5585 22958 5602
rect 23000 5585 23017 5602
rect 23142 5585 23159 5602
rect 23173 5571 23174 5617
rect 23187 5557 23188 5631
rect 23201 5585 23218 5602
rect 23260 5585 23277 5602
rect 23402 5585 23419 5602
rect 23433 5571 23434 5617
rect 23447 5557 23448 5631
rect 23461 5585 23478 5602
rect 23520 5585 23537 5602
rect 23662 5585 23679 5602
rect 23693 5571 23694 5617
rect 23707 5557 23708 5631
rect 23721 5585 23738 5602
rect 23780 5585 23797 5602
rect 23922 5585 23939 5602
rect 23953 5571 23954 5617
rect 23967 5557 23968 5631
rect 23981 5585 23998 5602
rect 24040 5585 24057 5602
rect 24182 5585 24199 5602
rect 24213 5571 24214 5617
rect 24227 5557 24228 5631
rect 24241 5585 24258 5602
rect 24300 5585 24317 5602
rect 24442 5585 24459 5602
rect 24473 5571 24474 5617
rect 24487 5557 24488 5631
rect 24501 5585 24518 5602
rect 24560 5585 24577 5602
rect 24702 5585 24719 5602
rect 24733 5571 24734 5617
rect 24747 5557 24748 5631
rect 24761 5585 24778 5602
rect 24820 5585 24837 5602
rect 24962 5585 24979 5602
rect 24993 5571 24994 5617
rect 25007 5557 25008 5631
rect 25021 5585 25038 5602
rect 25080 5585 25097 5602
rect 25222 5585 25239 5602
rect 25253 5571 25254 5617
rect 25267 5557 25268 5631
rect 25281 5585 25298 5602
rect 25340 5585 25357 5602
rect 25482 5585 25499 5602
rect 25513 5571 25514 5617
rect 25527 5557 25528 5631
rect 25541 5585 25558 5602
rect 25600 5585 25617 5602
rect 25742 5585 25759 5602
rect 25773 5571 25774 5617
rect 25787 5557 25788 5631
rect 25801 5585 25818 5602
rect 25860 5585 25877 5602
rect 26002 5585 26019 5602
rect 26033 5571 26034 5617
rect 26047 5557 26048 5631
rect 26061 5585 26078 5602
rect 26120 5585 26137 5602
rect 26262 5585 26279 5602
rect 26293 5571 26294 5617
rect 26307 5557 26308 5631
rect 26321 5585 26338 5602
rect 26380 5585 26397 5602
rect 26522 5585 26539 5602
rect 26553 5571 26554 5617
rect 26567 5557 26568 5631
rect 26581 5585 26598 5602
rect 26640 5585 26657 5602
rect 26782 5585 26799 5602
rect 26813 5571 26814 5617
rect 26827 5557 26828 5631
rect 26841 5585 26858 5602
rect 26900 5585 26917 5602
rect 27042 5585 27059 5602
rect 27073 5571 27074 5617
rect 27087 5557 27088 5631
rect 27101 5585 27118 5602
rect 27160 5585 27177 5602
rect 27302 5585 27319 5602
rect 27333 5571 27334 5617
rect 27347 5557 27348 5631
rect 27361 5585 27378 5602
rect 27420 5585 27437 5602
rect 27562 5585 27579 5602
rect 27593 5571 27594 5617
rect 27607 5557 27608 5631
rect 27621 5585 27638 5602
rect 27680 5585 27697 5602
rect 27822 5585 27839 5602
rect 27853 5571 27854 5617
rect 27867 5557 27868 5631
rect 27881 5585 27898 5602
rect 27940 5585 27957 5602
rect 28082 5585 28099 5602
rect 28113 5571 28114 5617
rect 28127 5557 28128 5631
rect 28141 5585 28158 5602
rect 28200 5585 28217 5602
rect 28342 5585 28359 5602
rect 28373 5571 28374 5617
rect 28387 5557 28388 5631
rect 28401 5585 28418 5602
rect 28460 5585 28477 5602
rect 28602 5585 28619 5602
rect 28633 5571 28634 5617
rect 28647 5557 28648 5631
rect 28661 5585 28678 5602
rect 28720 5585 28737 5602
rect 28862 5585 28879 5602
rect 28893 5571 28894 5617
rect 28907 5557 28908 5631
rect 28921 5585 28938 5602
rect 28980 5585 28997 5602
rect 29122 5585 29139 5602
rect 29153 5571 29154 5617
rect 29167 5557 29168 5631
rect 29181 5585 29198 5602
rect 29240 5585 29257 5602
rect 29382 5585 29399 5602
rect 29413 5571 29414 5617
rect 29427 5557 29428 5631
rect 29441 5585 29458 5602
rect 29500 5585 29517 5602
rect 29642 5585 29659 5602
rect 29673 5571 29674 5617
rect 29687 5557 29688 5631
rect 29701 5585 29718 5602
rect 29760 5585 29777 5602
rect 29902 5585 29919 5602
rect 29933 5571 29934 5617
rect 29947 5557 29948 5631
rect 29961 5585 29978 5602
rect 30020 5585 30037 5602
rect 30162 5585 30179 5602
rect 30193 5571 30194 5617
rect 30207 5557 30208 5631
rect 30221 5585 30238 5602
rect 30280 5585 30297 5602
rect 30422 5585 30439 5602
rect 30453 5571 30454 5617
rect 30467 5557 30468 5631
rect 30481 5585 30498 5602
rect 30540 5585 30557 5602
rect 30682 5585 30699 5602
rect 30713 5571 30714 5617
rect 30727 5557 30728 5631
rect 30741 5585 30758 5602
rect 30800 5585 30817 5602
rect 30942 5585 30959 5602
rect 30973 5571 30974 5617
rect 30987 5557 30988 5631
rect 31001 5585 31018 5602
rect 31060 5585 31077 5602
rect 31202 5585 31219 5602
rect 31233 5571 31234 5617
rect 31247 5557 31248 5631
rect 31261 5585 31278 5602
rect 31320 5585 31337 5602
rect 31462 5585 31479 5602
rect 31493 5571 31494 5617
rect 31507 5557 31508 5631
rect 31521 5585 31538 5602
rect 31580 5585 31597 5602
rect 1808 5541 1852 5542
rect 1808 5519 1809 5541
rect 1851 5519 1852 5541
rect 1281 5491 1298 5508
rect 1340 5491 1357 5508
rect 1595 5491 1612 5508
rect 1654 5491 1671 5508
rect 1909 5491 1926 5508
rect 1968 5491 1985 5508
rect 2223 5491 2240 5508
rect 2282 5491 2299 5508
rect 2537 5491 2554 5508
rect 2596 5491 2613 5508
rect 4283 5470 4300 5487
rect 4342 5470 4359 5487
rect 11987 5471 12004 5488
rect 12046 5471 12063 5488
rect 11523 5451 11540 5468
rect 11700 5451 11717 5468
rect 1379 5399 1434 5408
rect 1579 5390 1675 5408
rect 1693 5399 1748 5408
rect 1893 5390 1989 5408
rect 2007 5399 2062 5408
rect 2207 5390 2303 5408
rect 2321 5399 2376 5408
rect 2521 5390 2617 5408
rect 2635 5399 2690 5408
rect 11612 5396 11613 5411
rect 14867 5401 14868 5415
rect 15127 5401 15128 5415
rect 15387 5401 15388 5415
rect 15647 5401 15648 5415
rect 15907 5401 15908 5415
rect 16167 5401 16168 5415
rect 16427 5401 16428 5415
rect 16687 5401 16688 5415
rect 16947 5401 16948 5415
rect 17207 5401 17208 5415
rect 17467 5401 17468 5415
rect 17727 5401 17728 5415
rect 17987 5401 17988 5415
rect 18247 5401 18248 5415
rect 18507 5401 18508 5415
rect 18767 5401 18768 5415
rect 19027 5401 19028 5415
rect 19287 5401 19288 5415
rect 19547 5401 19548 5415
rect 19807 5401 19808 5415
rect 20067 5401 20068 5415
rect 20327 5401 20328 5415
rect 20587 5401 20588 5415
rect 20847 5401 20848 5415
rect 21107 5401 21108 5415
rect 21367 5401 21368 5415
rect 21627 5401 21628 5415
rect 21887 5401 21888 5415
rect 22147 5401 22148 5415
rect 22407 5401 22408 5415
rect 22667 5401 22668 5415
rect 22927 5401 22928 5415
rect 23187 5401 23188 5415
rect 23447 5401 23448 5415
rect 23707 5401 23708 5415
rect 23967 5401 23968 5415
rect 24227 5401 24228 5415
rect 24487 5401 24488 5415
rect 24747 5401 24748 5415
rect 25007 5401 25008 5415
rect 25267 5401 25268 5415
rect 25527 5401 25528 5415
rect 25787 5401 25788 5415
rect 26047 5401 26048 5415
rect 26307 5401 26308 5415
rect 26567 5401 26568 5415
rect 26827 5401 26828 5415
rect 27087 5401 27088 5415
rect 27347 5401 27348 5415
rect 27607 5401 27608 5415
rect 27867 5401 27868 5415
rect 28127 5401 28128 5415
rect 28387 5401 28388 5415
rect 28647 5401 28648 5415
rect 28907 5401 28908 5415
rect 29167 5401 29168 5415
rect 29427 5401 29428 5415
rect 29687 5401 29688 5415
rect 29947 5401 29948 5415
rect 30207 5401 30208 5415
rect 30467 5401 30468 5415
rect 30727 5401 30728 5415
rect 30987 5401 30988 5415
rect 31247 5401 31248 5415
rect 31507 5401 31508 5415
rect 12085 5379 12140 5388
rect 1357 5369 1366 5370
rect 1671 5369 1680 5370
rect 1985 5369 1994 5370
rect 2299 5369 2308 5370
rect 2613 5369 2622 5370
rect 14822 5369 14839 5386
rect 12047 5350 12063 5367
rect 14852 5355 14854 5401
rect 14866 5355 14868 5401
rect 14881 5369 14898 5386
rect 15082 5369 15099 5386
rect 15112 5355 15114 5401
rect 15126 5355 15128 5401
rect 15141 5369 15158 5386
rect 15342 5369 15359 5386
rect 15372 5355 15374 5401
rect 15386 5355 15388 5401
rect 15401 5369 15418 5386
rect 15602 5369 15619 5386
rect 15632 5355 15634 5401
rect 15646 5355 15648 5401
rect 15661 5369 15678 5386
rect 15862 5369 15879 5386
rect 15892 5355 15894 5401
rect 15906 5355 15908 5401
rect 15921 5369 15938 5386
rect 16122 5369 16139 5386
rect 16152 5355 16154 5401
rect 16166 5355 16168 5401
rect 16181 5369 16198 5386
rect 16382 5369 16399 5386
rect 16412 5355 16414 5401
rect 16426 5355 16428 5401
rect 16441 5369 16458 5386
rect 16642 5369 16659 5386
rect 16672 5355 16674 5401
rect 16686 5355 16688 5401
rect 16701 5369 16718 5386
rect 16902 5369 16919 5386
rect 16932 5355 16934 5401
rect 16946 5355 16948 5401
rect 16961 5369 16978 5386
rect 17162 5369 17179 5386
rect 17192 5355 17194 5401
rect 17206 5355 17208 5401
rect 17221 5369 17238 5386
rect 17422 5369 17439 5386
rect 17452 5355 17454 5401
rect 17466 5355 17468 5401
rect 17481 5369 17498 5386
rect 17682 5369 17699 5386
rect 17712 5355 17714 5401
rect 17726 5355 17728 5401
rect 17741 5369 17758 5386
rect 17942 5369 17959 5386
rect 17972 5355 17974 5401
rect 17986 5355 17988 5401
rect 18001 5369 18018 5386
rect 18202 5369 18219 5386
rect 18232 5355 18234 5401
rect 18246 5355 18248 5401
rect 18261 5369 18278 5386
rect 18462 5369 18479 5386
rect 18492 5355 18494 5401
rect 18506 5355 18508 5401
rect 18521 5369 18538 5386
rect 18722 5369 18739 5386
rect 18752 5355 18754 5401
rect 18766 5355 18768 5401
rect 18781 5369 18798 5386
rect 18982 5369 18999 5386
rect 19012 5355 19014 5401
rect 19026 5355 19028 5401
rect 19041 5369 19058 5386
rect 19242 5369 19259 5386
rect 19272 5355 19274 5401
rect 19286 5355 19288 5401
rect 19301 5369 19318 5386
rect 19502 5369 19519 5386
rect 19532 5355 19534 5401
rect 19546 5355 19548 5401
rect 19561 5369 19578 5386
rect 19762 5369 19779 5386
rect 19792 5355 19794 5401
rect 19806 5355 19808 5401
rect 19821 5369 19838 5386
rect 20022 5369 20039 5386
rect 20052 5355 20054 5401
rect 20066 5355 20068 5401
rect 20081 5369 20098 5386
rect 20282 5369 20299 5386
rect 20312 5355 20314 5401
rect 20326 5355 20328 5401
rect 20341 5369 20358 5386
rect 20542 5369 20559 5386
rect 20572 5355 20574 5401
rect 20586 5355 20588 5401
rect 20601 5369 20618 5386
rect 20802 5369 20819 5386
rect 20832 5355 20834 5401
rect 20846 5355 20848 5401
rect 20861 5369 20878 5386
rect 21062 5369 21079 5386
rect 21092 5355 21094 5401
rect 21106 5355 21108 5401
rect 21121 5369 21138 5386
rect 21322 5369 21339 5386
rect 21352 5355 21354 5401
rect 21366 5355 21368 5401
rect 21381 5369 21398 5386
rect 21582 5369 21599 5386
rect 21612 5355 21614 5401
rect 21626 5355 21628 5401
rect 21641 5369 21658 5386
rect 21842 5369 21859 5386
rect 21872 5355 21874 5401
rect 21886 5355 21888 5401
rect 21901 5369 21918 5386
rect 22102 5369 22119 5386
rect 22132 5355 22134 5401
rect 22146 5355 22148 5401
rect 22161 5369 22178 5386
rect 22362 5369 22379 5386
rect 22392 5355 22394 5401
rect 22406 5355 22408 5401
rect 22421 5369 22438 5386
rect 22622 5369 22639 5386
rect 22652 5355 22654 5401
rect 22666 5355 22668 5401
rect 22681 5369 22698 5386
rect 22882 5369 22899 5386
rect 22912 5355 22914 5401
rect 22926 5355 22928 5401
rect 22941 5369 22958 5386
rect 23142 5369 23159 5386
rect 23172 5355 23174 5401
rect 23186 5355 23188 5401
rect 23201 5369 23218 5386
rect 23402 5369 23419 5386
rect 23432 5355 23434 5401
rect 23446 5355 23448 5401
rect 23461 5369 23478 5386
rect 23662 5369 23679 5386
rect 23692 5355 23694 5401
rect 23706 5355 23708 5401
rect 23721 5369 23738 5386
rect 23922 5369 23939 5386
rect 23952 5355 23954 5401
rect 23966 5355 23968 5401
rect 23981 5369 23998 5386
rect 24182 5369 24199 5386
rect 24212 5355 24214 5401
rect 24226 5355 24228 5401
rect 24241 5369 24258 5386
rect 24442 5369 24459 5386
rect 24472 5355 24474 5401
rect 24486 5355 24488 5401
rect 24501 5369 24518 5386
rect 24702 5369 24719 5386
rect 24732 5355 24734 5401
rect 24746 5355 24748 5401
rect 24761 5369 24778 5386
rect 24962 5369 24979 5386
rect 24992 5355 24994 5401
rect 25006 5355 25008 5401
rect 25021 5369 25038 5386
rect 25222 5369 25239 5386
rect 25252 5355 25254 5401
rect 25266 5355 25268 5401
rect 25281 5369 25298 5386
rect 25482 5369 25499 5386
rect 25512 5355 25514 5401
rect 25526 5355 25528 5401
rect 25541 5369 25558 5386
rect 25742 5369 25759 5386
rect 25772 5355 25774 5401
rect 25786 5355 25788 5401
rect 25801 5369 25818 5386
rect 26002 5369 26019 5386
rect 26032 5355 26034 5401
rect 26046 5355 26048 5401
rect 26061 5369 26078 5386
rect 26262 5369 26279 5386
rect 26292 5355 26294 5401
rect 26306 5355 26308 5401
rect 26321 5369 26338 5386
rect 26522 5369 26539 5386
rect 26552 5355 26554 5401
rect 26566 5355 26568 5401
rect 26581 5369 26598 5386
rect 26782 5369 26799 5386
rect 26812 5355 26814 5401
rect 26826 5355 26828 5401
rect 26841 5369 26858 5386
rect 27042 5369 27059 5386
rect 27072 5355 27074 5401
rect 27086 5355 27088 5401
rect 27101 5369 27118 5386
rect 27302 5369 27319 5386
rect 27332 5355 27334 5401
rect 27346 5355 27348 5401
rect 27361 5369 27378 5386
rect 27562 5369 27579 5386
rect 27592 5355 27594 5401
rect 27606 5355 27608 5401
rect 27621 5369 27638 5386
rect 27822 5369 27839 5386
rect 27852 5355 27854 5401
rect 27866 5355 27868 5401
rect 27881 5369 27898 5386
rect 28082 5369 28099 5386
rect 28112 5355 28114 5401
rect 28126 5355 28128 5401
rect 28141 5369 28158 5386
rect 28342 5369 28359 5386
rect 28372 5355 28374 5401
rect 28386 5355 28388 5401
rect 28401 5369 28418 5386
rect 28602 5369 28619 5386
rect 28632 5355 28634 5401
rect 28646 5355 28648 5401
rect 28661 5369 28678 5386
rect 28862 5369 28879 5386
rect 28892 5355 28894 5401
rect 28906 5355 28908 5401
rect 28921 5369 28938 5386
rect 29122 5369 29139 5386
rect 29152 5355 29154 5401
rect 29166 5355 29168 5401
rect 29181 5369 29198 5386
rect 29382 5369 29399 5386
rect 29412 5355 29414 5401
rect 29426 5355 29428 5401
rect 29441 5369 29458 5386
rect 29642 5369 29659 5386
rect 29672 5355 29674 5401
rect 29686 5355 29688 5401
rect 29701 5369 29718 5386
rect 29902 5369 29919 5386
rect 29932 5355 29934 5401
rect 29946 5355 29948 5401
rect 29961 5369 29978 5386
rect 30162 5369 30179 5386
rect 30192 5355 30194 5401
rect 30206 5355 30208 5401
rect 30221 5369 30238 5386
rect 30422 5369 30439 5386
rect 30452 5355 30454 5401
rect 30466 5355 30468 5401
rect 30481 5369 30498 5386
rect 30682 5369 30699 5386
rect 30712 5355 30714 5401
rect 30726 5355 30728 5401
rect 30741 5369 30758 5386
rect 30942 5369 30959 5386
rect 30972 5355 30974 5401
rect 30986 5355 30988 5401
rect 31001 5369 31018 5386
rect 31202 5369 31219 5386
rect 31232 5355 31234 5401
rect 31246 5355 31248 5401
rect 31261 5369 31278 5386
rect 31462 5369 31479 5386
rect 31492 5355 31494 5401
rect 31506 5355 31508 5401
rect 31521 5369 31538 5386
rect 12047 5349 12080 5350
rect 4367 5347 4368 5348
rect 14867 5341 14868 5355
rect 15127 5341 15128 5355
rect 15387 5341 15388 5355
rect 15647 5341 15648 5355
rect 15907 5341 15908 5355
rect 16167 5341 16168 5355
rect 16427 5341 16428 5355
rect 16687 5341 16688 5355
rect 16947 5341 16948 5355
rect 17207 5341 17208 5355
rect 17467 5341 17468 5355
rect 17727 5341 17728 5355
rect 17987 5341 17988 5355
rect 18247 5341 18248 5355
rect 18507 5341 18508 5355
rect 18767 5341 18768 5355
rect 19027 5341 19028 5355
rect 19287 5341 19288 5355
rect 19547 5341 19548 5355
rect 19807 5341 19808 5355
rect 20067 5341 20068 5355
rect 20327 5341 20328 5355
rect 20587 5341 20588 5355
rect 20847 5341 20848 5355
rect 21107 5341 21108 5355
rect 21367 5341 21368 5355
rect 21627 5341 21628 5355
rect 21887 5341 21888 5355
rect 22147 5341 22148 5355
rect 22407 5341 22408 5355
rect 22667 5341 22668 5355
rect 22927 5341 22928 5355
rect 23187 5341 23188 5355
rect 23447 5341 23448 5355
rect 23707 5341 23708 5355
rect 23967 5341 23968 5355
rect 24227 5341 24228 5355
rect 24487 5341 24488 5355
rect 24747 5341 24748 5355
rect 25007 5341 25008 5355
rect 25267 5341 25268 5355
rect 25527 5341 25528 5355
rect 25787 5341 25788 5355
rect 26047 5341 26048 5355
rect 26307 5341 26308 5355
rect 26567 5341 26568 5355
rect 26827 5341 26828 5355
rect 27087 5341 27088 5355
rect 27347 5341 27348 5355
rect 27607 5341 27608 5355
rect 27867 5341 27868 5355
rect 28127 5341 28128 5355
rect 28387 5341 28388 5355
rect 28647 5341 28648 5355
rect 28907 5341 28908 5355
rect 29167 5341 29168 5355
rect 29427 5341 29428 5355
rect 29687 5341 29688 5355
rect 29947 5341 29948 5355
rect 30207 5341 30208 5355
rect 30467 5341 30468 5355
rect 30727 5341 30728 5355
rect 30987 5341 30988 5355
rect 31247 5341 31248 5355
rect 31507 5341 31508 5355
rect 14852 5315 14853 5330
rect 15112 5315 15113 5330
rect 15372 5315 15373 5330
rect 15632 5315 15633 5330
rect 15892 5315 15893 5330
rect 16152 5315 16153 5330
rect 16412 5315 16413 5330
rect 16672 5315 16673 5330
rect 16932 5315 16933 5330
rect 17192 5315 17193 5330
rect 17452 5315 17453 5330
rect 17712 5315 17713 5330
rect 17972 5315 17973 5330
rect 18232 5315 18233 5330
rect 18492 5315 18493 5330
rect 18752 5315 18753 5330
rect 19012 5315 19013 5330
rect 19272 5315 19273 5330
rect 19532 5315 19533 5330
rect 19792 5315 19793 5330
rect 20052 5315 20053 5330
rect 20312 5315 20313 5330
rect 20572 5315 20573 5330
rect 20832 5315 20833 5330
rect 21092 5315 21093 5330
rect 21352 5315 21353 5330
rect 21612 5315 21613 5330
rect 21872 5315 21873 5330
rect 22132 5315 22133 5330
rect 22392 5315 22393 5330
rect 22652 5315 22653 5330
rect 22912 5315 22913 5330
rect 23172 5315 23173 5330
rect 23432 5315 23433 5330
rect 23692 5315 23693 5330
rect 23952 5315 23953 5330
rect 24212 5315 24213 5330
rect 24472 5315 24473 5330
rect 24732 5315 24733 5330
rect 24992 5315 24993 5330
rect 25252 5315 25253 5330
rect 25512 5315 25513 5330
rect 25772 5315 25773 5330
rect 26032 5315 26033 5330
rect 26292 5315 26293 5330
rect 26552 5315 26553 5330
rect 26812 5315 26813 5330
rect 27072 5315 27073 5330
rect 27332 5315 27333 5330
rect 27592 5315 27593 5330
rect 27852 5315 27853 5330
rect 28112 5315 28113 5330
rect 28372 5315 28373 5330
rect 28632 5315 28633 5330
rect 28892 5315 28893 5330
rect 29152 5315 29153 5330
rect 29412 5315 29413 5330
rect 29672 5315 29673 5330
rect 29932 5315 29933 5330
rect 30192 5315 30193 5330
rect 30452 5315 30453 5330
rect 30712 5315 30713 5330
rect 30972 5315 30973 5330
rect 31232 5315 31233 5330
rect 31492 5315 31493 5330
rect 4381 5292 4436 5301
rect 11627 5270 11649 5285
rect 11627 5264 11628 5270
rect 11725 5251 11734 5252
rect 11675 5243 11700 5250
rect 11717 5243 11742 5250
rect 11675 5235 11742 5243
rect 11599 5234 11742 5235
rect 1281 5213 1298 5230
rect 1340 5213 1357 5230
rect 1595 5213 1612 5230
rect 1654 5213 1671 5230
rect 1909 5213 1926 5230
rect 1968 5213 1985 5230
rect 2223 5213 2240 5230
rect 2282 5213 2299 5230
rect 2537 5213 2554 5230
rect 2596 5213 2613 5230
rect 11676 5225 11725 5234
rect 11599 5217 11607 5218
rect 11633 5217 11666 5218
rect 10418 5213 10462 5214
rect 1644 5171 1645 5193
rect 1687 5171 1688 5193
rect 4283 5192 4300 5209
rect 4342 5192 4359 5209
rect 10418 5191 10419 5213
rect 10461 5191 10462 5213
rect 11320 5213 11364 5214
rect 11320 5191 11321 5213
rect 11363 5191 11364 5213
rect 11523 5193 11540 5210
rect 11582 5193 11599 5210
rect 11641 5193 11658 5210
rect 11687 5188 11725 5225
rect 11987 5193 12004 5210
rect 12046 5193 12063 5210
rect 11717 5180 11725 5188
rect 1644 5170 1688 5171
rect 1146 5155 1273 5156
rect 1306 5155 1390 5156
rect 1423 5155 1587 5156
rect 1620 5155 1704 5156
rect 1737 5155 1901 5156
rect 1934 5155 2018 5156
rect 2051 5155 2215 5156
rect 2248 5155 2332 5156
rect 2365 5155 2529 5156
rect 2562 5155 2646 5156
rect 2679 5155 2716 5156
rect 4148 5155 4275 5156
rect 4308 5155 4392 5156
rect 4425 5155 7259 5156
rect 4656 5085 4673 5102
rect 4715 5085 4732 5102
rect 4970 5085 4987 5102
rect 5039 5085 5056 5102
rect 5107 5085 5124 5102
rect 10362 5101 10414 5106
rect 11332 5101 11384 5106
rect 1179 5082 1187 5083
rect 1215 5082 1223 5083
rect 1179 5040 1180 5082
rect 1222 5040 1223 5082
rect 1281 5064 1298 5081
rect 1340 5064 1357 5081
rect 1595 5064 1612 5081
rect 1654 5064 1671 5081
rect 1909 5064 1926 5081
rect 1968 5064 1985 5081
rect 2223 5064 2240 5081
rect 2282 5064 2299 5081
rect 2537 5064 2554 5081
rect 2596 5064 2613 5081
rect 4283 5065 4300 5082
rect 4401 5065 4418 5082
rect 5362 5077 5379 5094
rect 5431 5077 5448 5094
rect 5509 5077 5526 5094
rect 5587 5077 5604 5094
rect 5665 5077 5682 5094
rect 5733 5077 5750 5094
rect 5988 5077 6005 5094
rect 6057 5077 6074 5094
rect 6135 5077 6152 5094
rect 6213 5077 6230 5094
rect 6291 5077 6308 5094
rect 6369 5077 6386 5094
rect 6447 5077 6464 5094
rect 6525 5077 6542 5094
rect 6603 5077 6620 5094
rect 6681 5077 6698 5094
rect 6759 5077 6776 5094
rect 6837 5077 6854 5094
rect 6915 5077 6932 5094
rect 6993 5077 7010 5094
rect 7071 5077 7088 5094
rect 7139 5077 7156 5094
rect 10332 5071 10444 5076
rect 11302 5071 11414 5076
rect 11717 5070 11725 5074
rect 5078 5052 5079 5067
rect 1179 5039 1223 5040
rect 4292 5031 4426 5036
rect 5704 5035 5705 5050
rect 7110 5035 7111 5050
rect 11523 5044 11540 5061
rect 11582 5044 11599 5061
rect 11641 5044 11658 5061
rect 11676 5046 11725 5070
rect 11599 5036 11607 5037
rect 11633 5036 11666 5037
rect 4372 5010 4373 5025
rect 11687 5020 11725 5046
rect 11987 5044 12004 5061
rect 12046 5044 12063 5061
rect 11599 5019 11751 5020
rect 4440 4993 4495 5002
rect 4640 4984 4736 5002
rect 4754 4993 4809 5002
rect 5032 4984 5050 5002
rect 5146 4993 5201 5002
rect 5772 4993 5827 5018
rect 7178 4993 7233 5018
rect 11675 5011 11742 5019
rect 11612 4990 11613 5005
rect 11627 4990 11628 5005
rect 11675 5004 11700 5011
rect 11717 5004 11742 5011
rect 1357 4941 1366 4942
rect 1671 4941 1680 4942
rect 1985 4941 1994 4942
rect 2299 4941 2308 4942
rect 2613 4941 2622 4942
rect 5719 4912 5720 4927
rect 7125 4912 7126 4927
rect 12047 4922 12063 4939
rect 12047 4921 12080 4922
rect 1379 4886 1434 4895
rect 1579 4886 1675 4904
rect 1693 4886 1748 4895
rect 1893 4886 1989 4904
rect 2007 4886 2062 4895
rect 2207 4886 2303 4904
rect 2321 4886 2376 4895
rect 2521 4886 2617 4904
rect 2635 4886 2690 4895
rect 4372 4878 4373 4880
rect 4387 4878 4388 4893
rect 5093 4878 5094 4893
rect 5431 4882 5583 4883
rect 5600 4882 5750 4883
rect 6057 4882 6599 4883
rect 6616 4882 7156 4883
rect 4427 4873 4435 4874
rect 4347 4857 4414 4864
rect 11627 4858 11628 4873
rect 12085 4866 12140 4875
rect 4344 4849 4417 4857
rect 4434 4856 4444 4857
rect 4347 4832 4413 4849
rect 4451 4839 4461 4857
rect 4352 4824 4413 4832
rect 4283 4807 4300 4824
rect 4342 4822 4418 4824
rect 4342 4807 4373 4822
rect 1281 4786 1298 4803
rect 1340 4786 1357 4803
rect 1595 4786 1612 4803
rect 1654 4786 1671 4803
rect 1909 4786 1926 4803
rect 1968 4786 1985 4803
rect 2223 4786 2240 4803
rect 2282 4786 2299 4803
rect 2537 4786 2554 4803
rect 2596 4786 2613 4803
rect 4352 4802 4373 4807
rect 4388 4807 4418 4822
rect 4656 4807 4673 4824
rect 4715 4807 4732 4824
rect 4970 4807 4987 4824
rect 5039 4807 5056 4824
rect 5107 4807 5124 4824
rect 5362 4823 5379 4840
rect 5431 4823 5448 4840
rect 5509 4823 5526 4840
rect 5587 4823 5604 4840
rect 5665 4823 5682 4840
rect 5733 4823 5750 4840
rect 5988 4823 6005 4840
rect 6057 4823 6074 4840
rect 6135 4823 6152 4840
rect 6213 4823 6230 4840
rect 6291 4823 6308 4840
rect 6369 4823 6386 4840
rect 6447 4823 6464 4840
rect 6525 4823 6542 4840
rect 6603 4823 6620 4840
rect 6681 4823 6698 4840
rect 6759 4823 6776 4840
rect 6837 4823 6854 4840
rect 6915 4823 6932 4840
rect 6993 4823 7010 4840
rect 7071 4823 7088 4840
rect 7139 4823 7156 4840
rect 4388 4802 4409 4807
rect 11523 4786 11540 4803
rect 11700 4786 11717 4803
rect 10254 4761 10255 4783
rect 10297 4761 10298 4783
rect 10254 4760 10298 4761
rect 11402 4761 11403 4783
rect 11445 4761 11446 4783
rect 11987 4766 12004 4783
rect 12046 4766 12063 4783
rect 11402 4760 11446 4761
rect 1146 4749 1273 4750
rect 1306 4749 1390 4750
rect 1423 4749 1587 4750
rect 1620 4749 1704 4750
rect 1737 4749 1901 4750
rect 1934 4749 2018 4750
rect 2051 4749 2215 4750
rect 2248 4749 2332 4750
rect 2365 4749 2529 4750
rect 2562 4749 2646 4750
rect 2679 4749 2716 4750
rect 4148 4749 4275 4750
rect 4308 4749 4393 4750
rect 4426 4749 4451 4750
rect 4484 4749 4648 4750
rect 4681 4749 4765 4750
rect 4798 4749 4962 4750
rect 4995 4749 5099 4750
rect 5132 4749 5157 4750
rect 5190 4749 5354 4750
rect 5387 4749 5501 4750
rect 5533 4749 5657 4750
rect 5689 4749 5783 4750
rect 5816 4749 5980 4750
rect 6013 4749 6127 4750
rect 6159 4749 6283 4750
rect 6315 4749 6439 4750
rect 6471 4749 6595 4750
rect 6627 4749 6751 4750
rect 6783 4749 6907 4750
rect 6939 4749 7063 4750
rect 7095 4749 7189 4750
rect 7222 4749 7259 4750
rect 15032 4740 15049 4757
rect 15091 4740 15108 4757
rect 15292 4740 15309 4757
rect 15351 4740 15368 4757
rect 15552 4740 15569 4757
rect 15611 4740 15628 4757
rect 15812 4740 15829 4757
rect 15871 4740 15888 4757
rect 16072 4740 16089 4757
rect 16131 4740 16148 4757
rect 16332 4740 16349 4757
rect 16391 4740 16408 4757
rect 16592 4740 16609 4757
rect 16651 4740 16668 4757
rect 16852 4740 16869 4757
rect 16911 4740 16928 4757
rect 17112 4740 17129 4757
rect 17171 4740 17188 4757
rect 17372 4740 17389 4757
rect 17431 4740 17448 4757
rect 17632 4740 17649 4757
rect 17691 4740 17708 4757
rect 17892 4740 17909 4757
rect 17951 4740 17968 4757
rect 18152 4740 18169 4757
rect 18211 4740 18228 4757
rect 18412 4740 18429 4757
rect 18471 4740 18488 4757
rect 18672 4740 18689 4757
rect 18731 4740 18748 4757
rect 18932 4740 18949 4757
rect 18991 4740 19008 4757
rect 19192 4740 19209 4757
rect 19251 4740 19268 4757
rect 19452 4740 19469 4757
rect 19511 4740 19528 4757
rect 19712 4740 19729 4757
rect 19771 4740 19788 4757
rect 19972 4740 19989 4757
rect 20031 4740 20048 4757
rect 20232 4740 20249 4757
rect 20291 4740 20308 4757
rect 20492 4740 20509 4757
rect 20551 4740 20568 4757
rect 20752 4740 20769 4757
rect 20811 4740 20828 4757
rect 21012 4740 21029 4757
rect 21071 4740 21088 4757
rect 21272 4740 21289 4757
rect 21331 4740 21348 4757
rect 21532 4740 21549 4757
rect 21591 4740 21608 4757
rect 21792 4740 21809 4757
rect 21851 4740 21868 4757
rect 22052 4740 22069 4757
rect 22111 4740 22128 4757
rect 22312 4740 22329 4757
rect 22371 4740 22388 4757
rect 22572 4740 22589 4757
rect 22631 4740 22648 4757
rect 22832 4740 22849 4757
rect 22891 4740 22908 4757
rect 23092 4740 23109 4757
rect 23151 4740 23168 4757
rect 23352 4740 23369 4757
rect 23411 4740 23428 4757
rect 23612 4740 23629 4757
rect 23671 4740 23688 4757
rect 23872 4740 23889 4757
rect 23931 4740 23948 4757
rect 24132 4740 24149 4757
rect 24191 4740 24208 4757
rect 24392 4740 24409 4757
rect 24451 4740 24468 4757
rect 24652 4740 24669 4757
rect 24711 4740 24728 4757
rect 24912 4740 24929 4757
rect 24971 4740 24988 4757
rect 25172 4740 25189 4757
rect 25231 4740 25248 4757
rect 25432 4740 25449 4757
rect 25491 4740 25508 4757
rect 25692 4740 25709 4757
rect 25751 4740 25768 4757
rect 25952 4740 25969 4757
rect 26011 4740 26028 4757
rect 26212 4740 26229 4757
rect 26271 4740 26288 4757
rect 26472 4740 26489 4757
rect 26531 4740 26548 4757
rect 26732 4740 26749 4757
rect 26791 4740 26808 4757
rect 26992 4740 27009 4757
rect 27051 4740 27068 4757
rect 27252 4740 27269 4757
rect 27311 4740 27328 4757
rect 27512 4740 27529 4757
rect 27571 4740 27588 4757
rect 27772 4740 27789 4757
rect 27831 4740 27848 4757
rect 28032 4740 28049 4757
rect 28091 4740 28108 4757
rect 28292 4740 28309 4757
rect 28351 4740 28368 4757
rect 28552 4740 28569 4757
rect 28611 4740 28628 4757
rect 28812 4740 28829 4757
rect 28871 4740 28888 4757
rect 29072 4740 29089 4757
rect 29131 4740 29148 4757
rect 29332 4740 29349 4757
rect 29391 4740 29408 4757
rect 29592 4740 29609 4757
rect 29651 4740 29668 4757
rect 29852 4740 29869 4757
rect 29911 4740 29928 4757
rect 30112 4740 30129 4757
rect 30171 4740 30188 4757
rect 30372 4740 30389 4757
rect 30431 4740 30448 4757
rect 30632 4740 30649 4757
rect 30691 4740 30708 4757
rect 30892 4740 30909 4757
rect 30951 4740 30968 4757
rect 31152 4740 31169 4757
rect 31211 4740 31228 4757
rect 31412 4740 31429 4757
rect 31471 4740 31488 4757
rect 10336 4721 10380 4722
rect 10336 4699 10337 4721
rect 10379 4699 10380 4721
rect 1281 4679 1298 4696
rect 1340 4679 1357 4696
rect 1595 4679 1612 4696
rect 1654 4679 1671 4696
rect 1909 4679 1926 4696
rect 1968 4679 1985 4696
rect 2223 4679 2240 4696
rect 2282 4679 2299 4696
rect 2537 4679 2554 4696
rect 2596 4679 2613 4696
rect 4477 4684 4485 4688
rect 4283 4658 4300 4675
rect 4342 4658 4359 4675
rect 4401 4658 4418 4675
rect 4436 4660 4485 4684
rect 4359 4650 4367 4651
rect 4393 4650 4426 4651
rect 4447 4634 4485 4660
rect 11987 4659 12004 4676
rect 12046 4659 12063 4676
rect 4747 4640 4764 4657
rect 4816 4640 4833 4657
rect 4894 4640 4911 4657
rect 4972 4640 4989 4657
rect 5050 4640 5067 4657
rect 5128 4640 5145 4657
rect 5206 4640 5223 4657
rect 5284 4640 5301 4657
rect 5362 4640 5379 4657
rect 5440 4640 5457 4657
rect 5518 4640 5535 4657
rect 5586 4640 5603 4657
rect 11523 4639 11540 4656
rect 11700 4639 11717 4656
rect 4359 4633 4511 4634
rect 4435 4625 4502 4633
rect 4372 4604 4373 4619
rect 4387 4604 4388 4619
rect 4435 4618 4460 4625
rect 4477 4618 4502 4625
rect 4833 4614 4972 4615
rect 4989 4614 5128 4615
rect 5145 4614 5284 4615
rect 5301 4614 5440 4615
rect 5457 4614 5586 4615
rect 1379 4587 1434 4596
rect 1579 4578 1675 4596
rect 1693 4587 1748 4596
rect 1893 4578 1989 4596
rect 2007 4587 2062 4596
rect 2207 4578 2303 4596
rect 2321 4587 2376 4596
rect 2521 4578 2617 4596
rect 2635 4587 2690 4596
rect 11612 4584 11613 4599
rect 5557 4566 5558 4581
rect 12085 4567 12140 4576
rect 1357 4557 1366 4558
rect 1671 4557 1680 4558
rect 1985 4557 1994 4558
rect 2299 4557 2308 4558
rect 2613 4557 2622 4558
rect 12047 4538 12063 4555
rect 12047 4537 12080 4538
rect 4387 4472 4388 4487
rect 5572 4462 5573 4464
rect 5625 4462 5680 4489
rect 4705 4460 5680 4462
rect 5572 4449 5573 4460
rect 11627 4458 11649 4473
rect 11627 4452 11628 4458
rect 11725 4439 11734 4440
rect 11675 4431 11700 4438
rect 11717 4431 11742 4438
rect 11675 4423 11742 4431
rect 11599 4422 11742 4423
rect 1281 4401 1298 4418
rect 1340 4401 1357 4418
rect 1595 4401 1612 4418
rect 1654 4401 1671 4418
rect 1909 4401 1926 4418
rect 1968 4401 1985 4418
rect 2223 4401 2240 4418
rect 2282 4401 2299 4418
rect 2537 4401 2554 4418
rect 2596 4401 2613 4418
rect 4283 4400 4300 4417
rect 4460 4400 4477 4417
rect 11676 4413 11725 4422
rect 4747 4389 4764 4406
rect 4816 4389 4833 4406
rect 4894 4389 4911 4406
rect 4972 4389 4989 4406
rect 5050 4389 5067 4406
rect 5128 4389 5145 4406
rect 5206 4389 5223 4406
rect 5284 4389 5301 4406
rect 5362 4389 5379 4406
rect 5440 4389 5457 4406
rect 5518 4389 5535 4406
rect 5586 4389 5603 4406
rect 11599 4405 11607 4406
rect 11633 4405 11666 4406
rect 11523 4381 11540 4398
rect 11582 4381 11599 4398
rect 11641 4381 11658 4398
rect 11687 4376 11725 4413
rect 11987 4381 12004 4398
rect 12046 4381 12063 4398
rect 15032 4377 15049 4394
rect 15091 4377 15108 4394
rect 15292 4377 15309 4394
rect 15351 4377 15368 4394
rect 15552 4377 15569 4394
rect 15611 4377 15628 4394
rect 15812 4377 15829 4394
rect 15871 4377 15888 4394
rect 16072 4377 16089 4394
rect 16131 4377 16148 4394
rect 16332 4377 16349 4394
rect 16391 4377 16408 4394
rect 16592 4377 16609 4394
rect 16651 4377 16668 4394
rect 16852 4377 16869 4394
rect 16911 4377 16928 4394
rect 17112 4377 17129 4394
rect 17171 4377 17188 4394
rect 17372 4377 17389 4394
rect 17431 4377 17448 4394
rect 17632 4377 17649 4394
rect 17691 4377 17708 4394
rect 17892 4377 17909 4394
rect 17951 4377 17968 4394
rect 18152 4377 18169 4394
rect 18211 4377 18228 4394
rect 18412 4377 18429 4394
rect 18471 4377 18488 4394
rect 18672 4377 18689 4394
rect 18731 4377 18748 4394
rect 18932 4377 18949 4394
rect 18991 4377 19008 4394
rect 19192 4377 19209 4394
rect 19251 4377 19268 4394
rect 19452 4377 19469 4394
rect 19511 4377 19528 4394
rect 19712 4377 19729 4394
rect 19771 4377 19788 4394
rect 19972 4377 19989 4394
rect 20031 4377 20048 4394
rect 20232 4377 20249 4394
rect 20291 4377 20308 4394
rect 20492 4377 20509 4394
rect 20551 4377 20568 4394
rect 20752 4377 20769 4394
rect 20811 4377 20828 4394
rect 21012 4377 21029 4394
rect 21071 4377 21088 4394
rect 21272 4377 21289 4394
rect 21331 4377 21348 4394
rect 21532 4377 21549 4394
rect 21591 4377 21608 4394
rect 21792 4377 21809 4394
rect 21851 4377 21868 4394
rect 22052 4377 22069 4394
rect 22111 4377 22128 4394
rect 22312 4377 22329 4394
rect 22371 4377 22388 4394
rect 22572 4377 22589 4394
rect 22631 4377 22648 4394
rect 22832 4377 22849 4394
rect 22891 4377 22908 4394
rect 23092 4377 23109 4394
rect 23151 4377 23168 4394
rect 23352 4377 23369 4394
rect 23411 4377 23428 4394
rect 23612 4377 23629 4394
rect 23671 4377 23688 4394
rect 23872 4377 23889 4394
rect 23931 4377 23948 4394
rect 24132 4377 24149 4394
rect 24191 4377 24208 4394
rect 24392 4377 24409 4394
rect 24451 4377 24468 4394
rect 24652 4377 24669 4394
rect 24711 4377 24728 4394
rect 24912 4377 24929 4394
rect 24971 4377 24988 4394
rect 25172 4377 25189 4394
rect 25231 4377 25248 4394
rect 25432 4377 25449 4394
rect 25491 4377 25508 4394
rect 25692 4377 25709 4394
rect 25751 4377 25768 4394
rect 25952 4377 25969 4394
rect 26011 4377 26028 4394
rect 26212 4377 26229 4394
rect 26271 4377 26288 4394
rect 26472 4377 26489 4394
rect 26531 4377 26548 4394
rect 26732 4377 26749 4394
rect 26791 4377 26808 4394
rect 26992 4377 27009 4394
rect 27051 4377 27068 4394
rect 27252 4377 27269 4394
rect 27311 4377 27328 4394
rect 27512 4377 27529 4394
rect 27571 4377 27588 4394
rect 27772 4377 27789 4394
rect 27831 4377 27848 4394
rect 28032 4377 28049 4394
rect 28091 4377 28108 4394
rect 28292 4377 28309 4394
rect 28351 4377 28368 4394
rect 28552 4377 28569 4394
rect 28611 4377 28628 4394
rect 28812 4377 28829 4394
rect 28871 4377 28888 4394
rect 29072 4377 29089 4394
rect 29131 4377 29148 4394
rect 29332 4377 29349 4394
rect 29391 4377 29408 4394
rect 29592 4377 29609 4394
rect 29651 4377 29668 4394
rect 29852 4377 29869 4394
rect 29911 4377 29928 4394
rect 30112 4377 30129 4394
rect 30171 4377 30188 4394
rect 30372 4377 30389 4394
rect 30431 4377 30448 4394
rect 30632 4377 30649 4394
rect 30691 4377 30708 4394
rect 30892 4377 30909 4394
rect 30951 4377 30968 4394
rect 31152 4377 31169 4394
rect 31211 4377 31228 4394
rect 31412 4377 31429 4394
rect 31471 4377 31488 4394
rect 1726 4351 1727 4373
rect 1769 4351 1770 4373
rect 11717 4368 11725 4376
rect 1726 4350 1770 4351
rect 1146 4343 1273 4344
rect 1306 4343 1390 4344
rect 1423 4343 1587 4344
rect 1620 4343 1704 4344
rect 1737 4343 1901 4344
rect 1934 4343 2018 4344
rect 2051 4343 2215 4344
rect 2248 4343 2332 4344
rect 2365 4343 2529 4344
rect 2562 4343 2646 4344
rect 2679 4343 2716 4344
rect 4148 4343 4275 4344
rect 4308 4343 4739 4344
rect 4772 4343 4886 4344
rect 4918 4343 5042 4344
rect 5074 4343 5198 4344
rect 5230 4343 5354 4344
rect 5386 4343 5510 4344
rect 5542 4343 5636 4344
rect 5669 4343 5706 4344
rect 4283 4253 4300 4270
rect 4460 4253 4477 4270
rect 4747 4267 4764 4284
rect 4816 4267 4833 4284
rect 4894 4267 4911 4284
rect 4972 4267 4989 4284
rect 5050 4267 5067 4284
rect 5128 4267 5145 4284
rect 5196 4267 5213 4284
rect 4886 4258 4918 4259
rect 5042 4258 5074 4259
rect 11717 4258 11725 4262
rect 5127 4242 5128 4250
rect 4869 4241 4935 4242
rect 5025 4241 5091 4242
rect 5167 4226 5168 4241
rect 11523 4232 11540 4249
rect 11582 4232 11599 4249
rect 11641 4232 11658 4249
rect 11676 4234 11725 4258
rect 11599 4224 11607 4225
rect 11633 4224 11666 4225
rect 4372 4198 4373 4213
rect 11687 4208 11725 4234
rect 11987 4232 12004 4249
rect 12046 4232 12063 4249
rect 11599 4207 11751 4208
rect 5235 4181 5290 4200
rect 11675 4199 11742 4207
rect 11612 4178 11613 4193
rect 11627 4178 11628 4193
rect 11675 4192 11700 4199
rect 11717 4192 11742 4199
rect 15062 4197 15063 4212
rect 15322 4197 15323 4212
rect 15582 4197 15583 4212
rect 15842 4197 15843 4212
rect 16102 4197 16103 4212
rect 16362 4197 16363 4212
rect 16622 4197 16623 4212
rect 16882 4197 16883 4212
rect 17142 4197 17143 4212
rect 17402 4197 17403 4212
rect 17662 4197 17663 4212
rect 17922 4197 17923 4212
rect 18182 4197 18183 4212
rect 18442 4197 18443 4212
rect 18702 4197 18703 4212
rect 18962 4197 18963 4212
rect 19222 4197 19223 4212
rect 19482 4197 19483 4212
rect 19742 4197 19743 4212
rect 20002 4197 20003 4212
rect 20262 4197 20263 4212
rect 20522 4197 20523 4212
rect 20782 4197 20783 4212
rect 21042 4197 21043 4212
rect 21302 4197 21303 4212
rect 21562 4197 21563 4212
rect 21822 4197 21823 4212
rect 22082 4197 22083 4212
rect 22342 4197 22343 4212
rect 22602 4197 22603 4212
rect 22862 4197 22863 4212
rect 23122 4197 23123 4212
rect 23382 4197 23383 4212
rect 23642 4197 23643 4212
rect 23902 4197 23903 4212
rect 24162 4197 24163 4212
rect 24422 4197 24423 4212
rect 24682 4197 24683 4212
rect 24942 4197 24943 4212
rect 25202 4197 25203 4212
rect 25462 4197 25463 4212
rect 25722 4197 25723 4212
rect 25982 4197 25983 4212
rect 26242 4197 26243 4212
rect 26502 4197 26503 4212
rect 26762 4197 26763 4212
rect 27022 4197 27023 4212
rect 27282 4197 27283 4212
rect 27542 4197 27543 4212
rect 27802 4197 27803 4212
rect 28062 4197 28063 4212
rect 28322 4197 28323 4212
rect 28582 4197 28583 4212
rect 28842 4197 28843 4212
rect 29102 4197 29103 4212
rect 29362 4197 29363 4212
rect 29622 4197 29623 4212
rect 29882 4197 29883 4212
rect 30142 4197 30143 4212
rect 30402 4197 30403 4212
rect 30662 4197 30663 4212
rect 30922 4197 30923 4212
rect 31182 4197 31183 4212
rect 31442 4197 31443 4212
rect 12047 4110 12063 4127
rect 12047 4109 12080 4110
rect 5182 4094 5183 4109
rect 4387 4072 4409 4087
rect 4387 4066 4388 4072
rect 5144 4059 5145 4067
rect 4485 4053 4494 4054
rect 4435 4045 4460 4052
rect 4477 4045 4502 4052
rect 4833 4050 4858 4051
rect 4869 4050 4936 4051
rect 4947 4050 4972 4051
rect 4989 4050 5014 4051
rect 5025 4050 5092 4051
rect 5103 4050 5128 4051
rect 11627 4046 11628 4061
rect 12085 4054 12140 4063
rect 4435 4037 4502 4045
rect 4359 4036 4502 4037
rect 4436 4027 4485 4036
rect 4833 4033 4841 4034
rect 4886 4033 4919 4034
rect 4964 4033 4972 4034
rect 4989 4033 4997 4034
rect 5042 4033 5075 4034
rect 5120 4033 5128 4034
rect 4359 4019 4367 4020
rect 4393 4019 4426 4020
rect 4283 3995 4300 4012
rect 4342 3995 4359 4012
rect 4401 3995 4418 4012
rect 4447 3990 4485 4027
rect 4747 4009 4764 4026
rect 4816 4009 4833 4026
rect 4894 4009 4911 4026
rect 4972 4009 4989 4026
rect 5050 4009 5067 4026
rect 5128 4009 5145 4026
rect 5196 4009 5213 4026
rect 4477 3982 4485 3990
rect 11523 3974 11540 3991
rect 11700 3974 11717 3991
rect 11402 3941 11403 3963
rect 11445 3941 11446 3963
rect 11987 3954 12004 3971
rect 12046 3954 12063 3971
rect 11402 3940 11446 3941
rect 4148 3937 4275 3938
rect 4308 3937 4393 3938
rect 4426 3937 4739 3938
rect 4772 3937 4886 3938
rect 4918 3937 5042 3938
rect 5074 3937 5188 3938
rect 5221 3937 5246 3938
rect 5279 3937 5491 3938
rect 11402 3901 11446 3902
rect 11402 3879 11403 3901
rect 11445 3879 11446 3901
rect 4348 3863 4413 3872
rect 4283 3846 4300 3863
rect 4342 3846 4418 3863
rect 4352 3838 4413 3846
rect 4347 3831 4413 3838
rect 4688 3832 4705 3849
rect 4757 3832 4774 3849
rect 4835 3832 4852 3849
rect 4913 3832 4930 3849
rect 4991 3832 5008 3849
rect 5069 3832 5086 3849
rect 5147 3832 5164 3849
rect 5225 3832 5242 3849
rect 5303 3832 5320 3849
rect 5371 3832 5388 3849
rect 11987 3847 12004 3864
rect 12046 3847 12063 3864
rect 4347 3823 4409 3831
rect 11523 3827 11540 3844
rect 11700 3827 11717 3844
rect 4774 3824 4782 3825
rect 4827 3824 4860 3825
rect 4905 3824 4913 3825
rect 4930 3824 4938 3825
rect 4983 3824 5016 3825
rect 5061 3824 5069 3825
rect 5086 3824 5094 3825
rect 5139 3824 5172 3825
rect 5217 3824 5225 3825
rect 5242 3824 5250 3825
rect 5295 3824 5328 3825
rect 5363 3824 5371 3825
rect 4347 3821 4373 3823
rect 4344 3814 4373 3821
rect 4388 3821 4409 3823
rect 4388 3814 4417 3821
rect 4344 3813 4417 3814
rect 4444 3813 4452 3814
rect 4347 3806 4414 3813
rect 4372 3792 4373 3806
rect 4452 3805 4453 3813
rect 4774 3807 4799 3808
rect 4810 3807 4877 3808
rect 4888 3807 4913 3808
rect 4930 3807 4955 3808
rect 4966 3807 5033 3808
rect 5044 3807 5069 3808
rect 5086 3807 5111 3808
rect 5122 3807 5189 3808
rect 5200 3807 5225 3808
rect 5242 3807 5267 3808
rect 5278 3807 5345 3808
rect 5346 3807 5371 3808
rect 5342 3764 5343 3779
rect 11612 3772 11613 3787
rect 12085 3755 12140 3764
rect 12047 3726 12063 3743
rect 12047 3725 12080 3726
rect 4387 3660 4388 3675
rect 5410 3658 5465 3677
rect 5357 3632 5358 3647
rect 11627 3646 11649 3661
rect 11627 3640 11628 3646
rect 11725 3627 11734 3628
rect 11675 3619 11700 3626
rect 11717 3619 11742 3626
rect 4810 3616 4876 3617
rect 4966 3616 5032 3617
rect 5122 3616 5188 3617
rect 5278 3616 5344 3617
rect 11675 3611 11742 3619
rect 11599 3610 11742 3611
rect 4283 3588 4300 3605
rect 4401 3588 4418 3605
rect 11676 3601 11725 3610
rect 4827 3599 4859 3600
rect 4983 3599 5015 3600
rect 5139 3599 5171 3600
rect 5295 3599 5327 3600
rect 11599 3593 11607 3594
rect 11633 3593 11666 3594
rect 4688 3574 4705 3591
rect 4757 3574 4774 3591
rect 4835 3574 4852 3591
rect 4913 3574 4930 3591
rect 4991 3574 5008 3591
rect 5069 3574 5086 3591
rect 5147 3574 5164 3591
rect 5225 3574 5242 3591
rect 5303 3574 5320 3591
rect 5371 3574 5388 3591
rect 11523 3569 11540 3586
rect 11582 3569 11599 3586
rect 11641 3569 11658 3586
rect 11687 3564 11725 3601
rect 11987 3569 12004 3586
rect 12046 3569 12063 3586
rect 11717 3556 11725 3564
rect 2692 3531 3554 3532
rect 4148 3531 4275 3532
rect 4308 3531 4680 3532
rect 4713 3531 4827 3532
rect 4859 3531 4983 3532
rect 5015 3531 5139 3532
rect 5171 3531 5295 3532
rect 5327 3531 5421 3532
rect 5454 3531 5805 3532
rect 10418 3531 10419 3553
rect 10461 3531 10462 3553
rect 10418 3530 10462 3531
rect 11320 3531 11321 3553
rect 11363 3531 11364 3553
rect 11320 3530 11364 3531
rect 2827 3461 2844 3478
rect 2896 3461 2913 3478
rect 2964 3461 2981 3478
rect 3219 3455 3236 3472
rect 3288 3455 3305 3472
rect 3366 3455 3383 3472
rect 3434 3455 3451 3472
rect 4283 3461 4300 3478
rect 4342 3461 4359 3478
rect 3358 3446 3390 3447
rect 2935 3428 2936 3443
rect 4597 3441 4614 3458
rect 4715 3441 4732 3458
rect 5002 3455 5019 3472
rect 5071 3455 5088 3472
rect 5149 3455 5166 3472
rect 5227 3455 5244 3472
rect 5305 3455 5322 3472
rect 5383 3455 5400 3472
rect 5461 3455 5478 3472
rect 5539 3455 5556 3472
rect 5617 3455 5634 3472
rect 5685 3455 5702 3472
rect 5141 3446 5173 3447
rect 5297 3446 5329 3447
rect 5453 3446 5485 3447
rect 5609 3446 5641 3447
rect 3341 3429 3407 3430
rect 5124 3429 5190 3430
rect 5280 3429 5346 3430
rect 5436 3429 5502 3430
rect 5592 3429 5658 3430
rect 3405 3414 3406 3429
rect 5656 3414 5657 3429
rect 10553 3420 10570 3437
rect 10612 3420 10629 3437
rect 3003 3369 3058 3378
rect 3473 3369 3528 3388
rect 4686 3386 4687 3401
rect 10966 3394 11004 3462
rect 11717 3446 11725 3450
rect 11523 3420 11540 3437
rect 11582 3420 11599 3437
rect 11641 3420 11658 3437
rect 11676 3422 11725 3446
rect 11599 3412 11607 3413
rect 11633 3412 11666 3413
rect 11687 3396 11725 3422
rect 11987 3420 12004 3437
rect 12046 3420 12063 3437
rect 11599 3395 11751 3396
rect 4381 3369 4436 3378
rect 5724 3369 5779 3388
rect 11675 3387 11742 3395
rect 11612 3366 11613 3381
rect 11627 3366 11628 3381
rect 11675 3380 11700 3387
rect 11717 3380 11742 3387
rect 10613 3298 10629 3315
rect 12047 3298 12063 3315
rect 10613 3297 10646 3298
rect 12047 3297 12080 3298
rect 3420 3282 3421 3297
rect 5671 3282 5672 3297
rect 15069 3282 15085 3293
rect 15099 3282 15115 3293
rect 17149 3282 17165 3293
rect 17179 3282 17195 3293
rect 19229 3282 19245 3293
rect 19259 3282 19275 3293
rect 21309 3282 21325 3293
rect 21339 3282 21355 3293
rect 23389 3282 23405 3293
rect 23419 3282 23435 3293
rect 25469 3282 25485 3293
rect 25499 3282 25515 3293
rect 27549 3282 27565 3293
rect 27579 3282 27595 3293
rect 29629 3282 29645 3293
rect 29659 3282 29675 3293
rect 2950 3254 2951 3269
rect 2827 3183 2844 3200
rect 2896 3183 2913 3200
rect 2964 3183 2981 3200
rect 3041 3173 3047 3253
rect 3058 3190 3064 3270
rect 4686 3254 4687 3256
rect 4701 3254 4702 3269
rect 15075 3268 15085 3279
rect 15099 3268 15108 3279
rect 17155 3268 17165 3279
rect 17179 3268 17188 3279
rect 19235 3268 19245 3279
rect 19259 3268 19268 3279
rect 21315 3268 21325 3279
rect 21339 3268 21348 3279
rect 23395 3268 23405 3279
rect 23419 3268 23428 3279
rect 25475 3268 25485 3279
rect 25499 3268 25508 3279
rect 27555 3268 27565 3279
rect 27579 3268 27588 3279
rect 29635 3268 29645 3279
rect 29659 3268 29668 3279
rect 4749 3250 4750 3258
rect 4741 3249 4749 3250
rect 10651 3242 10706 3251
rect 3305 3238 3330 3239
rect 3341 3238 3408 3239
rect 3409 3238 3434 3239
rect 4661 3233 4728 3240
rect 5088 3238 5113 3239
rect 5124 3238 5191 3239
rect 5202 3238 5227 3239
rect 5244 3238 5269 3239
rect 5280 3238 5347 3239
rect 5358 3238 5383 3239
rect 5400 3238 5425 3239
rect 5436 3238 5503 3239
rect 5514 3238 5539 3239
rect 5556 3238 5581 3239
rect 5592 3238 5659 3239
rect 5660 3238 5685 3239
rect 11627 3234 11628 3249
rect 12085 3242 12140 3251
rect 15666 3245 15710 3246
rect 4658 3225 4731 3233
rect 3305 3221 3313 3222
rect 3358 3221 3391 3222
rect 3426 3221 3434 3222
rect 4661 3217 4727 3225
rect 15666 3223 15667 3245
rect 15709 3223 15710 3245
rect 17716 3245 17760 3246
rect 17716 3223 17717 3245
rect 17759 3223 17760 3245
rect 19766 3245 19810 3246
rect 19766 3223 19767 3245
rect 19809 3223 19810 3245
rect 21898 3245 21942 3246
rect 21898 3223 21899 3245
rect 21941 3223 21942 3245
rect 23948 3245 23992 3246
rect 23948 3223 23949 3245
rect 23991 3223 23992 3245
rect 25998 3245 26042 3246
rect 25998 3223 25999 3245
rect 26041 3223 26042 3245
rect 28048 3245 28092 3246
rect 28048 3223 28049 3245
rect 28091 3223 28092 3245
rect 30180 3245 30224 3246
rect 30180 3223 30181 3245
rect 30223 3223 30224 3245
rect 5088 3221 5096 3222
rect 5141 3221 5174 3222
rect 5219 3221 5227 3222
rect 5244 3221 5252 3222
rect 5297 3221 5330 3222
rect 5375 3221 5383 3222
rect 5400 3221 5408 3222
rect 5453 3221 5486 3222
rect 5531 3221 5539 3222
rect 5556 3221 5564 3222
rect 5609 3221 5642 3222
rect 5677 3221 5685 3222
rect 3219 3197 3236 3214
rect 3288 3197 3305 3214
rect 3366 3197 3383 3214
rect 3434 3197 3451 3214
rect 4045 3200 4727 3217
rect 4045 3198 4732 3200
rect 4045 3192 4687 3198
rect 4283 3187 4300 3192
rect 4342 3187 4359 3192
rect 4597 3187 4614 3192
rect 4656 3187 4687 3192
rect 4045 3178 4687 3187
rect 4702 3183 4732 3198
rect 5002 3197 5019 3214
rect 5071 3197 5088 3214
rect 5149 3197 5166 3214
rect 5227 3197 5244 3214
rect 5305 3197 5322 3214
rect 5383 3197 5400 3214
rect 5461 3197 5478 3214
rect 5539 3197 5556 3214
rect 5617 3197 5634 3214
rect 5685 3197 5702 3214
rect 4702 3178 4723 3183
rect 4045 3162 4672 3178
rect 11523 3162 11540 3179
rect 11700 3162 11717 3179
rect 1021 3097 1059 3137
rect 1076 3108 1093 3126
rect 1150 3108 1167 3126
rect 1219 3108 1236 3126
rect 1298 3108 1315 3126
rect 1371 3108 1388 3126
rect 1526 3108 1543 3126
rect 1605 3108 1622 3126
rect 1684 3108 1701 3126
rect 1799 3108 1816 3126
rect 1878 3108 1895 3126
rect 1951 3108 1968 3126
rect 2130 3108 2147 3126
rect 2209 3108 2226 3126
rect 2692 3125 2819 3126
rect 2852 3125 2956 3126
rect 2989 3125 3014 3126
rect 3047 3125 3211 3126
rect 3244 3125 3358 3126
rect 3390 3125 3484 3126
rect 3517 3125 3554 3126
rect 4148 3125 4275 3126
rect 4308 3125 4392 3126
rect 4425 3125 4589 3126
rect 4622 3125 4707 3126
rect 4740 3125 4994 3126
rect 5027 3125 5141 3126
rect 5173 3125 5297 3126
rect 5329 3125 5453 3126
rect 5485 3125 5609 3126
rect 5641 3125 5735 3126
rect 5768 3125 8684 3126
rect 10500 3121 10501 3143
rect 10543 3121 10544 3143
rect 10553 3142 10570 3159
rect 10612 3142 10629 3159
rect 11987 3142 12004 3159
rect 12046 3142 12063 3159
rect 10500 3120 10544 3121
rect 2827 3034 2844 3051
rect 2896 3034 2913 3051
rect 2964 3034 2981 3051
rect 2935 2980 2936 2995
rect 3041 2981 3047 3061
rect 3058 2964 3064 3044
rect 3219 3020 3236 3037
rect 3288 3020 3305 3037
rect 3366 3020 3383 3037
rect 3434 3020 3451 3037
rect 4283 3034 4300 3051
rect 4342 3034 4359 3051
rect 4597 3034 4614 3051
rect 4656 3034 4673 3051
rect 4911 3034 4928 3051
rect 4970 3034 4987 3051
rect 5225 3020 5242 3037
rect 5294 3020 5311 3037
rect 5372 3020 5389 3037
rect 5440 3020 5457 3037
rect 5695 3020 5712 3037
rect 5764 3020 5781 3037
rect 5842 3020 5859 3037
rect 5920 3020 5937 3037
rect 5998 3020 6015 3037
rect 6076 3020 6093 3037
rect 6154 3020 6171 3037
rect 6232 3020 6249 3037
rect 6310 3020 6327 3037
rect 6378 3020 6395 3037
rect 10553 3035 10570 3052
rect 10612 3035 10629 3052
rect 11987 3035 12004 3052
rect 12046 3035 12063 3052
rect 15461 3048 15498 3060
rect 17541 3048 17578 3060
rect 19621 3048 19658 3060
rect 21701 3048 21738 3060
rect 23781 3048 23818 3060
rect 25861 3048 25898 3060
rect 27941 3048 27978 3060
rect 30021 3048 30058 3060
rect 15461 3033 15499 3048
rect 17541 3033 17579 3048
rect 19621 3033 19659 3048
rect 21701 3033 21739 3048
rect 23781 3033 23819 3048
rect 25861 3033 25899 3048
rect 27941 3033 27979 3048
rect 30021 3033 30059 3048
rect 6633 3014 6650 3031
rect 6702 3014 6719 3031
rect 6780 3014 6797 3031
rect 6858 3014 6875 3031
rect 6936 3014 6953 3031
rect 7014 3014 7031 3031
rect 7092 3014 7109 3031
rect 7170 3014 7187 3031
rect 7248 3014 7265 3031
rect 7326 3014 7343 3031
rect 7404 3014 7421 3031
rect 7482 3014 7499 3031
rect 7560 3014 7577 3031
rect 7638 3014 7655 3031
rect 7716 3014 7733 3031
rect 7794 3014 7811 3031
rect 7872 3014 7889 3031
rect 7950 3014 7967 3031
rect 8028 3014 8045 3031
rect 8106 3014 8123 3031
rect 8184 3014 8201 3031
rect 8262 3014 8279 3031
rect 8340 3014 8357 3031
rect 8418 3014 8435 3031
rect 8496 3014 8513 3031
rect 8564 3014 8581 3031
rect 11523 3015 11540 3032
rect 11700 3015 11717 3032
rect 15460 3022 15499 3033
rect 17540 3022 17579 3033
rect 19620 3022 19659 3033
rect 21700 3022 21739 3033
rect 23780 3022 23819 3033
rect 25860 3022 25899 3033
rect 27940 3022 27979 3033
rect 30020 3022 30059 3033
rect 3305 3012 3313 3013
rect 3358 3012 3391 3013
rect 3426 3012 3434 3013
rect 5311 3012 5319 3013
rect 5364 3012 5397 3013
rect 5432 3012 5440 3013
rect 5781 3012 5789 3013
rect 5834 3012 5867 3013
rect 5912 3012 5920 3013
rect 5937 3012 5945 3013
rect 5990 3012 6023 3013
rect 6068 3012 6076 3013
rect 6093 3012 6101 3013
rect 6146 3012 6179 3013
rect 6224 3012 6232 3013
rect 6249 3012 6257 3013
rect 6302 3012 6335 3013
rect 6370 3012 6378 3013
rect 6719 3006 6727 3007
rect 6772 3006 6805 3007
rect 6850 3006 6858 3007
rect 6875 3006 6883 3007
rect 6928 3006 6961 3007
rect 7006 3006 7014 3007
rect 7031 3006 7039 3007
rect 7084 3006 7117 3007
rect 7162 3006 7170 3007
rect 7187 3006 7195 3007
rect 7240 3006 7273 3007
rect 7318 3006 7326 3007
rect 7343 3006 7351 3007
rect 7396 3006 7429 3007
rect 7474 3006 7482 3007
rect 7499 3006 7507 3007
rect 7552 3006 7585 3007
rect 7630 3006 7638 3007
rect 7655 3006 7663 3007
rect 7708 3006 7741 3007
rect 7786 3006 7794 3007
rect 7811 3006 7819 3007
rect 7864 3006 7897 3007
rect 7942 3006 7950 3007
rect 7967 3006 7975 3007
rect 8020 3006 8053 3007
rect 8098 3006 8106 3007
rect 8123 3006 8131 3007
rect 8176 3006 8209 3007
rect 8254 3006 8262 3007
rect 8279 3006 8287 3007
rect 8332 3006 8365 3007
rect 8410 3006 8418 3007
rect 8435 3006 8443 3007
rect 8488 3006 8521 3007
rect 8556 3006 8564 3007
rect 15473 3000 15499 3022
rect 17553 3000 17579 3022
rect 19633 3000 19659 3022
rect 21713 3000 21739 3022
rect 23793 3000 23819 3022
rect 25873 3000 25899 3022
rect 27953 3000 27979 3022
rect 30033 3000 30059 3022
rect 15584 2999 15628 3000
rect 3305 2995 3330 2996
rect 3341 2995 3408 2996
rect 3409 2995 3434 2996
rect 5311 2995 5336 2996
rect 5347 2995 5414 2996
rect 5415 2995 5440 2996
rect 5781 2995 5806 2996
rect 5817 2995 5884 2996
rect 5895 2995 5920 2996
rect 5937 2995 5962 2996
rect 5973 2995 6040 2996
rect 6051 2995 6076 2996
rect 6093 2995 6118 2996
rect 6129 2995 6196 2996
rect 6207 2995 6232 2996
rect 6249 2995 6274 2996
rect 6285 2995 6352 2996
rect 6353 2995 6378 2996
rect 6719 2989 6744 2990
rect 6755 2989 6822 2990
rect 6833 2989 6858 2990
rect 6875 2989 6900 2990
rect 6911 2989 6978 2990
rect 6989 2989 7014 2990
rect 7031 2989 7056 2990
rect 7067 2989 7134 2990
rect 7145 2989 7170 2990
rect 7187 2989 7212 2990
rect 7223 2989 7290 2990
rect 7301 2989 7326 2990
rect 7343 2989 7368 2990
rect 7379 2989 7446 2990
rect 7457 2989 7482 2990
rect 7499 2989 7524 2990
rect 7535 2989 7602 2990
rect 7613 2989 7638 2990
rect 7655 2989 7680 2990
rect 7691 2989 7758 2990
rect 7769 2989 7794 2990
rect 7811 2989 7836 2990
rect 7847 2989 7914 2990
rect 7925 2989 7950 2990
rect 7967 2989 7992 2990
rect 8003 2989 8070 2990
rect 8081 2989 8106 2990
rect 8123 2989 8148 2990
rect 8159 2989 8226 2990
rect 8237 2989 8262 2990
rect 8279 2989 8304 2990
rect 8315 2989 8382 2990
rect 8393 2989 8418 2990
rect 8435 2989 8460 2990
rect 8471 2989 8538 2990
rect 8539 2989 8564 2990
rect 15489 2983 15498 2999
rect 15584 2977 15585 2999
rect 15627 2977 15628 2999
rect 17470 2999 17514 3000
rect 19684 2999 19728 3000
rect 21734 2999 21778 3000
rect 17470 2977 17471 2999
rect 17513 2977 17514 2999
rect 17569 2983 17578 2999
rect 19649 2983 19658 2999
rect 19684 2977 19685 2999
rect 19727 2977 19728 2999
rect 21729 2983 21738 2999
rect 21734 2977 21735 2983
rect 21777 2977 21778 2999
rect 23784 2999 23828 3000
rect 25916 2999 25960 3000
rect 23784 2977 23785 2999
rect 23809 2983 23818 2999
rect 23827 2977 23828 2999
rect 25889 2983 25898 2999
rect 25916 2977 25917 2999
rect 25959 2977 25960 2999
rect 27884 2999 27928 3000
rect 27884 2977 27885 2999
rect 27927 2977 27928 2999
rect 27969 2983 27978 2999
rect 30049 2983 30058 2999
rect 3405 2952 3406 2967
rect 5411 2952 5412 2967
rect 6349 2952 6350 2967
rect 11612 2960 11613 2975
rect 8535 2940 8536 2955
rect 10651 2943 10706 2952
rect 12085 2943 12140 2952
rect 4186 2917 4230 2918
rect 4186 2895 4187 2917
rect 4229 2895 4230 2917
rect 10613 2914 10629 2931
rect 12047 2914 12063 2931
rect 14919 2923 14936 2932
rect 15083 2923 15100 2932
rect 16999 2923 17016 2932
rect 17163 2923 17180 2932
rect 19079 2923 19096 2932
rect 19243 2923 19260 2932
rect 21159 2923 21176 2932
rect 21323 2923 21340 2932
rect 23239 2923 23256 2932
rect 23403 2923 23420 2932
rect 25319 2923 25336 2932
rect 25483 2923 25500 2932
rect 27399 2923 27416 2932
rect 27563 2923 27580 2932
rect 29479 2923 29496 2932
rect 29643 2923 29660 2932
rect 10613 2913 10646 2914
rect 12047 2913 12080 2914
rect 14908 2885 14946 2923
rect 15073 2885 15111 2923
rect 16988 2885 17026 2923
rect 17153 2885 17191 2923
rect 19068 2885 19106 2923
rect 19233 2885 19271 2923
rect 21148 2885 21186 2923
rect 21313 2885 21351 2923
rect 23228 2885 23266 2923
rect 23393 2885 23431 2923
rect 25308 2885 25346 2923
rect 25473 2885 25511 2923
rect 27388 2885 27426 2923
rect 27553 2885 27591 2923
rect 29468 2885 29506 2923
rect 29633 2885 29671 2923
rect 14914 2878 14940 2885
rect 15079 2878 15105 2885
rect 16994 2878 17020 2885
rect 17159 2878 17185 2885
rect 19074 2878 19100 2885
rect 19239 2878 19265 2885
rect 21154 2878 21180 2885
rect 21319 2878 21345 2885
rect 23234 2878 23260 2885
rect 23399 2878 23425 2885
rect 25314 2878 25340 2885
rect 25479 2878 25505 2885
rect 27394 2878 27420 2885
rect 27559 2878 27585 2885
rect 29474 2878 29500 2885
rect 29639 2878 29665 2885
rect 3003 2856 3058 2865
rect 3473 2846 3528 2865
rect 4381 2856 4436 2865
rect 4581 2856 4677 2874
rect 4695 2856 4750 2865
rect 4895 2856 4991 2874
rect 5009 2856 5064 2865
rect 5479 2846 5534 2865
rect 6417 2846 6472 2865
rect 8550 2839 8551 2841
rect 8603 2839 8658 2865
rect 2950 2806 2951 2821
rect 3420 2820 3421 2835
rect 5426 2820 5427 2835
rect 6364 2820 6365 2835
rect 6591 2834 8658 2839
rect 11627 2834 11649 2849
rect 8550 2826 8551 2834
rect 11627 2828 11628 2834
rect 6702 2824 7634 2825
rect 7651 2824 8581 2825
rect 11725 2815 11734 2816
rect 11675 2807 11700 2814
rect 11717 2807 11742 2814
rect 3341 2804 3407 2805
rect 5347 2804 5413 2805
rect 5817 2804 5883 2805
rect 5973 2804 6039 2805
rect 6129 2804 6195 2805
rect 6285 2804 6351 2805
rect 11675 2799 11742 2807
rect 11599 2798 11742 2799
rect 11676 2789 11725 2798
rect 3358 2787 3390 2788
rect 5364 2787 5396 2788
rect 5834 2787 5866 2788
rect 5990 2787 6022 2788
rect 6146 2787 6178 2788
rect 6302 2787 6334 2788
rect 2827 2756 2844 2773
rect 2896 2756 2913 2773
rect 2964 2756 2981 2773
rect 3219 2762 3236 2779
rect 3288 2762 3305 2779
rect 3366 2762 3383 2779
rect 3434 2762 3451 2779
rect 4283 2756 4300 2773
rect 4342 2756 4359 2773
rect 4597 2756 4614 2773
rect 4656 2756 4673 2773
rect 4911 2756 4928 2773
rect 4970 2756 4987 2773
rect 5225 2762 5242 2779
rect 5294 2762 5311 2779
rect 5372 2762 5389 2779
rect 5440 2762 5457 2779
rect 5695 2762 5712 2779
rect 5764 2762 5781 2779
rect 5842 2762 5859 2779
rect 5920 2762 5937 2779
rect 5998 2762 6015 2779
rect 6076 2762 6093 2779
rect 6154 2762 6171 2779
rect 6232 2762 6249 2779
rect 6310 2762 6327 2779
rect 6378 2762 6395 2779
rect 6633 2766 6650 2783
rect 6702 2766 6719 2783
rect 6780 2766 6797 2783
rect 6858 2766 6875 2783
rect 6936 2766 6953 2783
rect 7014 2766 7031 2783
rect 7092 2766 7109 2783
rect 7170 2766 7187 2783
rect 7248 2766 7265 2783
rect 7326 2766 7343 2783
rect 7404 2766 7421 2783
rect 7482 2766 7499 2783
rect 7560 2766 7577 2783
rect 7638 2766 7655 2783
rect 7716 2766 7733 2783
rect 7794 2766 7811 2783
rect 7872 2766 7889 2783
rect 7950 2766 7967 2783
rect 8028 2766 8045 2783
rect 8106 2766 8123 2783
rect 8184 2766 8201 2783
rect 8262 2766 8279 2783
rect 8340 2766 8357 2783
rect 8418 2766 8435 2783
rect 8496 2766 8513 2783
rect 8564 2766 8581 2783
rect 11599 2781 11607 2782
rect 11633 2781 11666 2782
rect 10553 2757 10570 2774
rect 10612 2757 10629 2774
rect 11523 2757 11540 2774
rect 11582 2757 11599 2774
rect 11641 2757 11658 2774
rect 11687 2752 11725 2789
rect 11987 2757 12004 2774
rect 12046 2757 12063 2774
rect 3421 2745 3462 2746
rect 11717 2744 11725 2752
rect 15502 2753 15546 2754
rect 1070 2711 1071 2733
rect 1113 2711 1114 2733
rect 3407 2731 3448 2732
rect 2692 2719 2819 2720
rect 2852 2719 2956 2720
rect 2989 2719 3014 2720
rect 3047 2719 3211 2720
rect 3244 2719 3358 2720
rect 3390 2719 3484 2720
rect 3517 2719 3554 2720
rect 4148 2719 4275 2720
rect 4308 2719 4392 2720
rect 4425 2719 4589 2720
rect 4622 2719 4706 2720
rect 4739 2719 4903 2720
rect 4936 2719 5020 2720
rect 5053 2719 5217 2720
rect 5250 2719 5364 2720
rect 5396 2719 5490 2720
rect 5523 2719 5687 2720
rect 5720 2719 5834 2720
rect 5866 2719 5990 2720
rect 6022 2719 6146 2720
rect 6178 2719 6302 2720
rect 6334 2719 6428 2720
rect 6461 2719 6625 2720
rect 6658 2719 6772 2720
rect 6804 2719 6928 2720
rect 6960 2719 7084 2720
rect 7116 2719 7240 2720
rect 7272 2719 7396 2720
rect 7428 2719 7552 2720
rect 7584 2719 7708 2720
rect 7740 2719 7864 2720
rect 7896 2719 8020 2720
rect 8052 2719 8176 2720
rect 8208 2719 8332 2720
rect 8364 2719 8488 2720
rect 8520 2719 8614 2720
rect 8647 2719 8684 2720
rect 1070 2710 1114 2711
rect 10336 2711 10337 2733
rect 10379 2711 10380 2733
rect 10336 2710 10380 2711
rect 11320 2711 11321 2733
rect 11363 2711 11364 2733
rect 15502 2731 15503 2753
rect 15545 2731 15546 2753
rect 17798 2753 17842 2754
rect 17798 2731 17799 2753
rect 17841 2731 17842 2753
rect 19848 2753 19892 2754
rect 19848 2731 19849 2753
rect 19891 2731 19892 2753
rect 21570 2753 21614 2754
rect 21570 2731 21571 2753
rect 21613 2731 21614 2753
rect 24030 2753 24074 2754
rect 24030 2731 24031 2753
rect 24073 2731 24074 2753
rect 26080 2753 26124 2754
rect 26080 2731 26081 2753
rect 26123 2731 26124 2753
rect 28130 2753 28174 2754
rect 28130 2731 28131 2753
rect 28173 2731 28174 2753
rect 30262 2753 30306 2754
rect 30262 2731 30263 2753
rect 30305 2731 30306 2753
rect 11320 2710 11364 2711
rect 10418 2671 10462 2672
rect 10418 2649 10419 2671
rect 10461 2649 10462 2671
rect 11717 2634 11725 2638
rect 10553 2608 10570 2625
rect 10612 2608 10629 2625
rect 11523 2608 11540 2625
rect 11582 2608 11599 2625
rect 11641 2608 11658 2625
rect 11676 2610 11725 2634
rect 23456 2629 23457 2651
rect 23499 2629 23500 2651
rect 23456 2628 23500 2629
rect 25588 2629 25589 2651
rect 25631 2629 25632 2651
rect 25588 2628 25632 2629
rect 27638 2629 27639 2651
rect 27681 2629 27682 2651
rect 27638 2628 27682 2629
rect 29688 2629 29689 2651
rect 29731 2629 29732 2651
rect 29688 2628 29732 2629
rect 11599 2600 11607 2601
rect 11633 2600 11666 2601
rect 11687 2584 11725 2610
rect 11987 2608 12004 2625
rect 12046 2608 12063 2625
rect 16240 2589 16284 2590
rect 11599 2583 11751 2584
rect 11675 2575 11742 2583
rect 11612 2554 11613 2569
rect 11627 2554 11628 2569
rect 11675 2568 11700 2575
rect 11717 2568 11742 2575
rect 16240 2567 16241 2589
rect 16283 2567 16284 2589
rect 22062 2589 22106 2590
rect 22062 2567 22063 2589
rect 22105 2567 22106 2589
rect 10613 2486 10629 2503
rect 12047 2486 12063 2503
rect 10613 2485 10646 2486
rect 12047 2485 12080 2486
rect 10651 2430 10706 2439
rect 11627 2422 11628 2437
rect 12085 2430 12140 2439
rect 11523 2350 11540 2367
rect 11700 2350 11717 2367
rect 10553 2330 10570 2347
rect 10612 2330 10629 2347
rect 11987 2330 12004 2347
rect 12046 2330 12063 2347
rect 10254 2301 10255 2323
rect 10297 2301 10298 2323
rect 10254 2300 10298 2301
rect 11402 2301 11403 2323
rect 11445 2301 11446 2323
rect 15394 2314 15461 2317
rect 17474 2314 17541 2317
rect 19554 2314 19621 2317
rect 21634 2314 21701 2317
rect 23714 2314 23781 2317
rect 25794 2314 25861 2317
rect 27874 2314 27941 2317
rect 29954 2314 30021 2317
rect 15200 2309 15264 2314
rect 15394 2309 15573 2314
rect 15200 2304 15573 2309
rect 17280 2309 17344 2314
rect 17474 2309 17653 2314
rect 17280 2304 17653 2309
rect 19360 2309 19424 2314
rect 19554 2309 19733 2314
rect 19360 2304 19733 2309
rect 21440 2309 21504 2314
rect 21634 2309 21813 2314
rect 21440 2304 21813 2309
rect 23520 2309 23584 2314
rect 23714 2309 23893 2314
rect 23520 2304 23893 2309
rect 25600 2309 25664 2314
rect 25794 2309 25973 2314
rect 25600 2304 25973 2309
rect 27680 2309 27744 2314
rect 27874 2309 28053 2314
rect 27680 2304 28053 2309
rect 29760 2309 29824 2314
rect 29954 2309 30133 2314
rect 29760 2304 30133 2309
rect 11402 2300 11446 2301
rect 15411 2297 15444 2300
rect 17491 2297 17524 2300
rect 19571 2297 19604 2300
rect 21651 2297 21684 2300
rect 23731 2297 23764 2300
rect 25811 2297 25844 2300
rect 27891 2297 27924 2300
rect 29971 2297 30004 2300
rect 15217 2292 15247 2297
rect 15411 2292 15573 2297
rect 15217 2287 15573 2292
rect 17297 2292 17327 2297
rect 17491 2292 17653 2297
rect 17297 2287 17653 2292
rect 19377 2292 19407 2297
rect 19571 2292 19733 2297
rect 19377 2287 19733 2292
rect 21457 2292 21487 2297
rect 21651 2292 21813 2297
rect 21457 2287 21813 2292
rect 23537 2292 23567 2297
rect 23731 2292 23893 2297
rect 23537 2287 23893 2292
rect 25617 2292 25647 2297
rect 25811 2292 25973 2297
rect 25617 2287 25973 2292
rect 27697 2292 27727 2297
rect 27891 2292 28053 2297
rect 27697 2287 28053 2292
rect 29777 2292 29807 2297
rect 29971 2292 30133 2297
rect 29777 2287 30133 2292
rect 10500 2261 10544 2262
rect 10500 2239 10501 2261
rect 10543 2239 10544 2261
rect 15075 2236 15092 2239
rect 17155 2236 17172 2239
rect 19235 2236 19252 2239
rect 21315 2236 21332 2239
rect 23395 2236 23412 2239
rect 25475 2236 25492 2239
rect 27555 2236 27572 2239
rect 29635 2236 29652 2239
rect 15062 2235 15106 2236
rect 15062 2193 15063 2235
rect 15075 2206 15092 2235
rect 15105 2193 15106 2235
rect 15062 2192 15070 2193
rect 15098 2192 15106 2193
rect 17142 2235 17186 2236
rect 17142 2193 17143 2235
rect 17155 2206 17172 2235
rect 17185 2193 17186 2235
rect 17142 2192 17150 2193
rect 17178 2192 17186 2193
rect 19222 2235 19266 2236
rect 19222 2193 19223 2235
rect 19235 2206 19252 2235
rect 19265 2193 19266 2235
rect 19222 2192 19230 2193
rect 19258 2192 19266 2193
rect 21302 2235 21346 2236
rect 21302 2193 21303 2235
rect 21315 2206 21332 2235
rect 21345 2193 21346 2235
rect 21302 2192 21310 2193
rect 21338 2192 21346 2193
rect 23382 2235 23426 2236
rect 23382 2193 23383 2235
rect 23395 2206 23412 2235
rect 23425 2193 23426 2235
rect 23382 2192 23390 2193
rect 23418 2192 23426 2193
rect 25462 2235 25506 2236
rect 25462 2193 25463 2235
rect 25475 2206 25492 2235
rect 25505 2193 25506 2235
rect 25462 2192 25470 2193
rect 25498 2192 25506 2193
rect 27542 2235 27586 2236
rect 27542 2193 27543 2235
rect 27555 2206 27572 2235
rect 27585 2193 27586 2235
rect 27542 2192 27550 2193
rect 27578 2192 27586 2193
rect 29622 2235 29666 2236
rect 29622 2193 29623 2235
rect 29635 2206 29652 2235
rect 29665 2193 29666 2235
rect 29622 2192 29630 2193
rect 29658 2192 29666 2193
rect 23538 2055 23539 2077
rect 23581 2055 23582 2077
rect 23538 2054 23582 2055
rect 29770 2055 29771 2077
rect 29813 2055 29814 2077
rect 29770 2054 29814 2055
rect 21980 2015 22024 2016
rect 21980 1993 21981 2015
rect 22023 1993 22024 2015
rect 25998 2015 26042 2016
rect 25998 1993 25999 2015
rect 26041 1993 26042 2015
rect 28130 2015 28174 2016
rect 28130 1993 28131 2015
rect 28173 1993 28174 2015
rect 17806 1851 17850 1852
rect 17806 1809 17807 1851
rect 17849 1809 17850 1851
rect 17806 1808 17814 1809
rect 17842 1808 17850 1809
rect 21302 1851 21310 1852
rect 21338 1851 21346 1852
rect 21302 1809 21303 1851
rect 21345 1809 21346 1851
rect 21302 1808 21346 1809
rect 22466 1851 22510 1852
rect 22466 1809 22467 1851
rect 22509 1809 22510 1851
rect 22466 1808 22474 1809
rect 22502 1808 22510 1809
rect 29622 1851 29630 1852
rect 29658 1851 29666 1852
rect 29622 1809 29623 1851
rect 29665 1809 29666 1851
rect 29622 1808 29666 1809
rect 21301 1769 21345 1770
rect 21301 1727 21302 1769
rect 21344 1727 21345 1769
rect 21301 1726 21309 1727
rect 21337 1726 21345 1727
rect 27542 1769 27550 1770
rect 27578 1769 27586 1770
rect 27542 1727 27543 1769
rect 27585 1727 27586 1769
rect 27542 1726 27586 1727
rect 16641 1687 16685 1688
rect 16641 1645 16642 1687
rect 16684 1645 16685 1687
rect 16641 1644 16649 1645
rect 16677 1644 16685 1645
rect 19222 1687 19230 1688
rect 19258 1687 19266 1688
rect 19222 1645 19223 1687
rect 19265 1645 19266 1687
rect 19222 1644 19266 1645
rect 20136 1687 20180 1688
rect 20136 1645 20137 1687
rect 20179 1645 20180 1687
rect 20136 1644 20144 1645
rect 20172 1644 20180 1645
rect 25462 1687 25470 1688
rect 25498 1687 25506 1688
rect 25462 1645 25463 1687
rect 25505 1645 25506 1687
rect 25462 1644 25506 1645
rect 14311 1605 14355 1606
rect 14311 1563 14312 1605
rect 14354 1563 14355 1605
rect 14311 1562 14319 1563
rect 14347 1562 14355 1563
rect 15062 1605 15070 1606
rect 15098 1605 15106 1606
rect 15062 1563 15063 1605
rect 15105 1563 15106 1605
rect 15062 1562 15106 1563
rect 15476 1605 15520 1606
rect 15476 1563 15477 1605
rect 15519 1563 15520 1605
rect 15476 1562 15484 1563
rect 15512 1562 15520 1563
rect 17142 1605 17150 1606
rect 17178 1605 17186 1606
rect 17142 1563 17143 1605
rect 17185 1563 17186 1605
rect 17142 1562 17186 1563
rect 18971 1605 19015 1606
rect 18971 1563 18972 1605
rect 19014 1563 19015 1605
rect 18971 1562 18979 1563
rect 19007 1562 19015 1563
rect 23382 1605 23390 1606
rect 23418 1605 23426 1606
rect 23382 1563 23383 1605
rect 23425 1563 23426 1605
rect 23382 1562 23426 1563
rect 17716 1481 17717 1503
rect 17759 1481 17760 1503
rect 17716 1480 17760 1481
rect 19766 1481 19767 1503
rect 19809 1481 19810 1503
rect 19766 1480 19810 1481
rect 11010 1412 11012 1429
rect 12175 1412 12177 1429
rect 13340 1412 13342 1429
rect 14505 1412 14507 1429
rect 15670 1412 15672 1429
rect 16835 1412 16837 1429
rect 18000 1412 18002 1429
rect 19165 1412 19167 1429
rect 20330 1412 20332 1429
rect 21495 1412 21497 1429
rect 9926 1359 9970 1360
rect 9926 1337 9927 1359
rect 9969 1337 9970 1359
rect 10418 1359 10462 1360
rect 10418 1337 10419 1359
rect 10461 1337 10462 1359
rect 11000 1348 11002 1365
rect 10977 1315 10985 1348
rect 10994 1315 11002 1348
rect 11038 1346 11043 1373
rect 11156 1359 11200 1360
rect 11046 1346 11060 1348
rect 11007 1323 11022 1346
rect 11035 1323 11036 1340
rect 11038 1323 11060 1346
rect 9923 1235 9975 1253
rect 11038 1229 11043 1323
rect 11046 1298 11060 1323
rect 11063 1315 11077 1348
rect 11156 1337 11157 1359
rect 11199 1337 11200 1359
rect 11566 1359 11610 1360
rect 11566 1337 11567 1359
rect 11609 1337 11610 1359
rect 12165 1348 12167 1365
rect 12142 1315 12150 1348
rect 12159 1315 12167 1348
rect 12203 1346 12208 1373
rect 12304 1359 12348 1360
rect 12211 1346 12225 1348
rect 12172 1323 12187 1346
rect 12200 1323 12201 1340
rect 12203 1323 12225 1346
rect 11053 1223 11060 1298
rect 11070 1223 11077 1315
rect 11088 1235 11140 1253
rect 12203 1229 12208 1323
rect 12211 1298 12225 1323
rect 12228 1315 12242 1348
rect 12304 1337 12305 1359
rect 12347 1337 12348 1359
rect 12714 1359 12758 1360
rect 12714 1337 12715 1359
rect 12757 1337 12758 1359
rect 13330 1348 13332 1365
rect 13307 1315 13315 1348
rect 13324 1315 13332 1348
rect 13368 1346 13373 1373
rect 13452 1359 13496 1360
rect 13376 1346 13390 1348
rect 13337 1323 13352 1346
rect 13365 1323 13366 1340
rect 13368 1323 13390 1346
rect 12218 1223 12225 1298
rect 12235 1223 12242 1315
rect 12253 1235 12305 1253
rect 13368 1229 13373 1323
rect 13376 1298 13390 1323
rect 13393 1315 13407 1348
rect 13452 1337 13453 1359
rect 13495 1337 13496 1359
rect 13862 1359 13906 1360
rect 13862 1337 13863 1359
rect 13905 1337 13906 1359
rect 14495 1348 14497 1365
rect 14472 1315 14480 1348
rect 14489 1315 14497 1348
rect 14533 1346 14538 1373
rect 14600 1359 14644 1360
rect 14541 1346 14555 1348
rect 14502 1323 14517 1346
rect 14530 1323 14531 1340
rect 14533 1323 14555 1346
rect 13383 1223 13390 1298
rect 13400 1223 13407 1315
rect 14311 1267 14319 1268
rect 14347 1267 14355 1268
rect 13418 1235 13470 1253
rect 14311 1225 14312 1267
rect 14354 1225 14355 1267
rect 14533 1229 14538 1323
rect 14541 1298 14555 1323
rect 14558 1315 14572 1348
rect 14600 1337 14601 1359
rect 14643 1337 14644 1359
rect 15010 1359 15054 1360
rect 15010 1337 15011 1359
rect 15053 1337 15054 1359
rect 15660 1348 15662 1365
rect 15637 1315 15645 1348
rect 15654 1315 15662 1348
rect 15698 1346 15703 1373
rect 15748 1359 15792 1360
rect 15706 1346 15720 1348
rect 15667 1323 15682 1346
rect 15695 1323 15696 1340
rect 15698 1323 15720 1346
rect 14311 1224 14355 1225
rect 14548 1223 14555 1298
rect 14565 1223 14572 1315
rect 15476 1267 15484 1268
rect 15512 1267 15520 1268
rect 14583 1235 14635 1253
rect 15476 1225 15477 1267
rect 15519 1225 15520 1267
rect 15698 1229 15703 1323
rect 15706 1298 15720 1323
rect 15723 1315 15737 1348
rect 15748 1337 15749 1359
rect 15791 1337 15792 1359
rect 16240 1359 16284 1360
rect 16240 1337 16241 1359
rect 16283 1337 16284 1359
rect 16825 1348 16827 1365
rect 16802 1315 16810 1348
rect 16819 1315 16827 1348
rect 16863 1346 16868 1373
rect 16978 1359 17022 1360
rect 16871 1346 16885 1348
rect 16832 1323 16847 1346
rect 16860 1323 16861 1340
rect 16863 1323 16885 1346
rect 15476 1224 15520 1225
rect 15713 1223 15720 1298
rect 15730 1223 15737 1315
rect 16641 1267 16649 1268
rect 16677 1267 16685 1268
rect 15748 1235 15800 1253
rect 16641 1225 16642 1267
rect 16684 1225 16685 1267
rect 16863 1229 16868 1323
rect 16871 1298 16885 1323
rect 16888 1315 16902 1348
rect 16978 1337 16979 1359
rect 17021 1337 17022 1359
rect 17306 1359 17350 1360
rect 17306 1337 17307 1359
rect 17349 1337 17350 1359
rect 17990 1348 17992 1365
rect 17967 1315 17975 1348
rect 17984 1315 17992 1348
rect 18028 1346 18033 1373
rect 18044 1359 18088 1360
rect 18044 1348 18045 1359
rect 18036 1346 18050 1348
rect 17997 1323 18012 1346
rect 18025 1323 18026 1340
rect 18028 1323 18050 1346
rect 16641 1224 16685 1225
rect 16878 1223 16885 1298
rect 16895 1223 16902 1315
rect 17806 1267 17814 1268
rect 17842 1267 17850 1268
rect 16913 1235 16965 1253
rect 17806 1225 17807 1267
rect 17849 1225 17850 1267
rect 18028 1229 18033 1323
rect 18036 1298 18050 1323
rect 18053 1315 18067 1348
rect 18087 1337 18088 1359
rect 18536 1359 18580 1360
rect 18536 1337 18537 1359
rect 18579 1337 18580 1359
rect 19155 1348 19157 1365
rect 19132 1315 19140 1348
rect 19149 1315 19157 1348
rect 19193 1346 19198 1373
rect 19274 1359 19318 1360
rect 19201 1346 19215 1348
rect 19162 1323 19177 1346
rect 19190 1323 19191 1340
rect 19193 1323 19215 1346
rect 17806 1224 17850 1225
rect 18043 1223 18050 1298
rect 18060 1223 18067 1315
rect 18971 1267 18979 1268
rect 19007 1267 19015 1268
rect 18078 1235 18130 1253
rect 18971 1225 18972 1267
rect 19014 1225 19015 1267
rect 19193 1229 19198 1323
rect 19201 1298 19215 1323
rect 19218 1315 19232 1348
rect 19274 1337 19275 1359
rect 19317 1337 19318 1359
rect 19766 1359 19810 1360
rect 19766 1337 19767 1359
rect 19809 1337 19810 1359
rect 20320 1348 20322 1365
rect 20297 1315 20305 1348
rect 20314 1315 20322 1348
rect 20358 1346 20363 1373
rect 20422 1359 20466 1360
rect 20366 1346 20380 1348
rect 20327 1323 20342 1346
rect 20355 1323 20356 1340
rect 20358 1323 20380 1346
rect 18971 1224 19015 1225
rect 19208 1223 19215 1298
rect 19225 1223 19232 1315
rect 20136 1267 20144 1268
rect 20172 1267 20180 1268
rect 19243 1235 19295 1253
rect 20136 1225 20137 1267
rect 20179 1225 20180 1267
rect 20358 1229 20363 1323
rect 20366 1298 20380 1323
rect 20383 1315 20397 1348
rect 20422 1337 20423 1359
rect 20465 1337 20466 1359
rect 20914 1359 20958 1360
rect 20914 1337 20915 1359
rect 20957 1337 20958 1359
rect 21485 1348 21487 1365
rect 21462 1315 21470 1348
rect 21479 1315 21487 1348
rect 21523 1346 21528 1373
rect 21570 1359 21614 1360
rect 21531 1346 21545 1348
rect 21492 1323 21507 1346
rect 21520 1323 21521 1340
rect 21523 1323 21545 1346
rect 20136 1224 20180 1225
rect 20373 1223 20380 1298
rect 20390 1223 20397 1315
rect 21301 1267 21309 1268
rect 21337 1267 21345 1268
rect 20408 1235 20460 1253
rect 21301 1225 21302 1267
rect 21344 1225 21345 1267
rect 21523 1229 21528 1323
rect 21531 1298 21545 1323
rect 21548 1315 21562 1348
rect 21570 1337 21571 1359
rect 21613 1337 21614 1359
rect 22144 1359 22188 1360
rect 22144 1337 22145 1359
rect 22187 1337 22188 1359
rect 21301 1224 21345 1225
rect 21538 1223 21545 1298
rect 21555 1223 21562 1315
rect 22466 1267 22474 1268
rect 22502 1267 22510 1268
rect 21573 1235 21625 1253
rect 22466 1225 22467 1267
rect 22509 1225 22510 1267
rect 22466 1224 22510 1225
rect 9893 1205 10005 1223
rect 10982 1176 11015 1179
rect 10982 1163 11036 1176
rect 10988 1159 11022 1162
rect 10968 1149 11022 1159
rect 10989 1146 11022 1149
rect 10977 1058 10985 1108
rect 10994 1075 11002 1108
rect 11038 1106 11043 1214
rect 11053 1205 11170 1223
rect 11053 1197 11060 1205
rect 11052 1134 11060 1197
rect 11070 1180 11077 1205
rect 11069 1151 11077 1180
rect 12147 1176 12180 1179
rect 12147 1163 12201 1176
rect 12153 1159 12187 1162
rect 11053 1125 11060 1134
rect 11046 1106 11060 1125
rect 11070 1108 11077 1151
rect 12133 1149 12187 1159
rect 12154 1146 12187 1149
rect 11007 1083 11022 1106
rect 11035 1083 11036 1100
rect 11038 1083 11060 1106
rect 10500 1031 10544 1032
rect 10500 1009 10501 1031
rect 10543 1009 10544 1031
rect 10983 1028 10985 1058
rect 11000 1028 11002 1075
rect 11038 1054 11043 1083
rect 11046 1075 11060 1083
rect 11063 1075 11077 1108
rect 12142 1058 12150 1108
rect 12159 1075 12167 1108
rect 12203 1106 12208 1214
rect 12218 1205 12335 1223
rect 12218 1197 12225 1205
rect 12217 1134 12225 1197
rect 12235 1180 12242 1205
rect 12234 1151 12242 1180
rect 13312 1176 13345 1179
rect 13312 1163 13366 1176
rect 13318 1159 13352 1162
rect 12218 1125 12225 1134
rect 12211 1106 12225 1125
rect 12235 1108 12242 1151
rect 13298 1149 13352 1159
rect 13319 1146 13352 1149
rect 12172 1083 12187 1106
rect 12200 1083 12201 1100
rect 12203 1083 12225 1106
rect 11648 1031 11692 1032
rect 10989 1003 11005 1020
rect 11031 1003 11048 1020
rect 11049 1003 11066 1020
rect 11648 1009 11649 1031
rect 11691 1009 11692 1031
rect 12148 1028 12150 1058
rect 12165 1028 12167 1075
rect 12203 1054 12208 1083
rect 12211 1075 12225 1083
rect 12228 1075 12242 1108
rect 13307 1058 13315 1108
rect 13324 1075 13332 1108
rect 13368 1106 13373 1214
rect 13383 1205 13500 1223
rect 13383 1197 13390 1205
rect 13382 1134 13390 1197
rect 13400 1180 13407 1205
rect 13399 1151 13407 1180
rect 14477 1176 14510 1179
rect 14477 1163 14531 1176
rect 14483 1159 14517 1162
rect 13383 1125 13390 1134
rect 13376 1106 13390 1125
rect 13400 1108 13407 1151
rect 14463 1149 14517 1159
rect 14484 1146 14517 1149
rect 13337 1083 13352 1106
rect 13365 1083 13366 1100
rect 13368 1083 13390 1106
rect 12796 1031 12840 1032
rect 12154 1003 12170 1020
rect 12196 1003 12213 1020
rect 12214 1003 12231 1020
rect 12796 1009 12797 1031
rect 12839 1009 12840 1031
rect 13313 1028 13315 1058
rect 13330 1028 13332 1075
rect 13368 1054 13373 1083
rect 13376 1075 13390 1083
rect 13393 1075 13407 1108
rect 14472 1058 14480 1108
rect 14489 1075 14497 1108
rect 14533 1106 14538 1214
rect 14548 1205 14665 1223
rect 14548 1197 14555 1205
rect 14547 1134 14555 1197
rect 14565 1180 14572 1205
rect 14564 1151 14572 1180
rect 15642 1176 15675 1179
rect 15642 1163 15696 1176
rect 15648 1159 15682 1162
rect 14548 1125 14555 1134
rect 14541 1106 14555 1125
rect 14565 1108 14572 1151
rect 15628 1149 15682 1159
rect 15649 1146 15682 1149
rect 14502 1083 14517 1106
rect 14530 1083 14531 1100
rect 14533 1083 14555 1106
rect 13944 1031 13988 1032
rect 13319 1003 13335 1020
rect 13361 1003 13378 1020
rect 13379 1003 13396 1020
rect 13944 1009 13945 1031
rect 13987 1009 13988 1031
rect 14478 1028 14480 1058
rect 14495 1028 14497 1075
rect 14533 1054 14538 1083
rect 14541 1075 14555 1083
rect 14558 1075 14572 1108
rect 15637 1058 15645 1108
rect 15654 1075 15662 1108
rect 15698 1106 15703 1214
rect 15713 1205 15830 1223
rect 15713 1197 15720 1205
rect 15712 1134 15720 1197
rect 15730 1180 15737 1205
rect 15729 1151 15737 1180
rect 16807 1176 16840 1179
rect 16807 1163 16861 1176
rect 16813 1159 16847 1162
rect 15713 1125 15720 1134
rect 15706 1106 15720 1125
rect 15730 1108 15737 1151
rect 16793 1149 16847 1159
rect 16814 1146 16847 1149
rect 15667 1093 15682 1106
rect 15092 1031 15136 1032
rect 14484 1003 14500 1020
rect 14526 1003 14543 1020
rect 14544 1003 14561 1020
rect 15092 1009 15093 1031
rect 15135 1009 15136 1031
rect 15643 1028 15645 1058
rect 15660 1028 15662 1075
rect 15666 1083 15682 1093
rect 15695 1083 15696 1100
rect 15698 1083 15720 1106
rect 15666 1071 15667 1083
rect 15698 1071 15703 1083
rect 15706 1075 15720 1083
rect 15723 1075 15737 1108
rect 15709 1071 15710 1075
rect 15666 1070 15710 1071
rect 15698 1054 15703 1070
rect 16802 1058 16810 1108
rect 16819 1075 16827 1108
rect 16863 1106 16868 1214
rect 16878 1205 16995 1223
rect 16878 1197 16885 1205
rect 16877 1134 16885 1197
rect 16895 1180 16902 1205
rect 16894 1151 16902 1180
rect 17972 1176 18005 1179
rect 17972 1163 18026 1176
rect 17978 1159 18012 1162
rect 16878 1125 16885 1134
rect 16871 1106 16885 1125
rect 16895 1108 16902 1151
rect 17958 1149 18012 1159
rect 17979 1146 18012 1149
rect 16832 1083 16847 1106
rect 16860 1083 16861 1100
rect 16863 1083 16885 1106
rect 16322 1031 16366 1032
rect 15649 1003 15665 1020
rect 15691 1003 15708 1020
rect 15709 1003 15726 1020
rect 16322 1009 16323 1031
rect 16365 1009 16366 1031
rect 16808 1028 16810 1058
rect 16825 1028 16827 1075
rect 16863 1054 16868 1083
rect 16871 1075 16885 1083
rect 16888 1075 16902 1108
rect 17634 1071 17635 1093
rect 17677 1071 17678 1093
rect 17634 1070 17678 1071
rect 17967 1058 17975 1108
rect 17984 1075 17992 1108
rect 18028 1106 18033 1214
rect 18043 1205 18160 1223
rect 18043 1197 18050 1205
rect 18042 1134 18050 1197
rect 18060 1180 18067 1205
rect 18059 1151 18067 1180
rect 19137 1176 19170 1179
rect 19137 1163 19191 1176
rect 19143 1159 19177 1162
rect 18043 1125 18050 1134
rect 18036 1106 18050 1125
rect 18060 1108 18067 1151
rect 19123 1149 19177 1159
rect 19144 1146 19177 1149
rect 17997 1083 18012 1106
rect 18025 1083 18026 1100
rect 18028 1083 18050 1106
rect 17634 1031 17678 1032
rect 16814 1003 16830 1020
rect 16856 1003 16873 1020
rect 16874 1003 16891 1020
rect 17634 1009 17635 1031
rect 17677 1009 17678 1031
rect 17973 1028 17975 1058
rect 17990 1028 17992 1075
rect 18028 1054 18033 1083
rect 18036 1075 18050 1083
rect 18053 1075 18067 1108
rect 19132 1058 19140 1108
rect 19149 1075 19157 1108
rect 19193 1106 19198 1214
rect 19208 1205 19325 1223
rect 19208 1197 19215 1205
rect 19207 1134 19215 1197
rect 19225 1180 19232 1205
rect 19224 1151 19232 1180
rect 20302 1176 20335 1179
rect 20302 1163 20356 1176
rect 20308 1159 20342 1162
rect 19208 1125 19215 1134
rect 19201 1106 19215 1125
rect 19225 1108 19232 1151
rect 20288 1149 20342 1159
rect 20309 1146 20342 1149
rect 19162 1083 19177 1106
rect 19190 1083 19191 1100
rect 19193 1083 19215 1106
rect 18618 1031 18662 1032
rect 17979 1003 17995 1020
rect 18021 1003 18038 1020
rect 18039 1003 18056 1020
rect 18618 1009 18619 1031
rect 18661 1009 18662 1031
rect 19138 1028 19140 1058
rect 19155 1028 19157 1075
rect 19193 1054 19198 1083
rect 19201 1075 19215 1083
rect 19218 1075 19232 1108
rect 19848 1071 19849 1093
rect 19891 1071 19892 1093
rect 19848 1070 19892 1071
rect 20297 1058 20305 1108
rect 20314 1075 20322 1108
rect 20358 1106 20363 1214
rect 20373 1205 20490 1223
rect 20373 1197 20380 1205
rect 20372 1134 20380 1197
rect 20390 1180 20397 1205
rect 20389 1151 20397 1180
rect 21467 1176 21500 1179
rect 21467 1163 21521 1176
rect 21473 1159 21507 1162
rect 20373 1125 20380 1134
rect 20366 1106 20380 1125
rect 20390 1108 20397 1151
rect 21453 1149 21507 1159
rect 21474 1146 21507 1149
rect 20327 1083 20342 1106
rect 20355 1083 20356 1100
rect 20358 1083 20380 1106
rect 19602 1031 19646 1032
rect 19144 1003 19160 1020
rect 19186 1003 19203 1020
rect 19204 1003 19221 1020
rect 19602 1009 19603 1031
rect 19645 1009 19646 1031
rect 20303 1028 20305 1058
rect 20320 1028 20322 1075
rect 20358 1054 20363 1083
rect 20366 1075 20380 1083
rect 20383 1075 20397 1108
rect 21462 1058 21470 1108
rect 21479 1075 21487 1108
rect 21523 1106 21528 1214
rect 21538 1205 21655 1223
rect 21538 1197 21545 1205
rect 21537 1134 21545 1197
rect 21555 1180 21562 1205
rect 21554 1151 21562 1180
rect 21538 1125 21545 1134
rect 21531 1106 21545 1125
rect 21555 1108 21562 1151
rect 21492 1083 21507 1106
rect 21520 1083 21521 1100
rect 21523 1083 21545 1106
rect 20832 1031 20876 1032
rect 20309 1003 20325 1020
rect 20351 1003 20368 1020
rect 20369 1003 20386 1020
rect 20832 1009 20833 1031
rect 20875 1009 20876 1031
rect 21468 1028 21470 1058
rect 21485 1028 21487 1075
rect 21523 1054 21528 1083
rect 21531 1075 21545 1083
rect 21548 1075 21562 1108
rect 22062 1031 22106 1032
rect 21474 1003 21490 1020
rect 21516 1003 21533 1020
rect 21534 1003 21551 1020
rect 22062 1009 22063 1031
rect 22105 1009 22106 1031
<< metal2 >>
rect 8809 2905 8823 14379
rect 8898 10622 8912 14401
rect 8964 10622 8978 14781
rect 9030 10622 9044 15213
rect 9096 10622 9110 15593
rect 9162 10622 9176 16025
rect 12938 5771 12952 6907
rect 13920 4958 13934 6048
rect 14002 4146 14016 6048
rect 14084 4523 14098 6048
rect 8750 2891 8823 2905
rect 8809 1208 8823 2891
<< metal3 >>
rect 164 24518 32852 24734
rect 574 24108 32442 24324
rect 14514 23832 14648 23914
rect 14760 23832 14894 23914
rect 15006 23862 15632 23914
rect 15006 23832 15140 23862
rect 14048 23780 15140 23832
rect 15252 23780 15386 23862
rect 15498 23832 15632 23862
rect 15744 23832 15878 23914
rect 15498 23780 15878 23832
rect 16072 23862 16452 23914
rect 16072 23780 16206 23862
rect 16318 23832 16452 23862
rect 16564 23862 17190 23914
rect 16564 23832 16698 23862
rect 16318 23780 16698 23832
rect 16810 23780 16944 23862
rect 17056 23832 17190 23862
rect 17302 23832 17518 23914
rect 17630 23862 18010 23914
rect 17630 23832 17764 23862
rect 17056 23780 17764 23832
rect 17876 23832 18010 23862
rect 18122 23832 18256 23914
rect 18368 23862 18748 23914
rect 18368 23832 18502 23862
rect 17876 23780 18502 23832
rect 18614 23832 18748 23862
rect 18942 23862 19322 23914
rect 18942 23832 19076 23862
rect 18614 23780 19076 23832
rect 19188 23832 19322 23862
rect 19434 23832 19568 23914
rect 19680 23832 19814 23914
rect 19926 23832 20060 23914
rect 20172 23832 20306 23914
rect 19188 23780 20306 23832
rect 20500 23832 20634 23914
rect 20746 23832 20880 23914
rect 20992 23832 21126 23914
rect 21238 23862 21618 23914
rect 21238 23832 21372 23862
rect 20500 23780 21372 23832
rect 21484 23832 21618 23862
rect 21730 23832 21864 23914
rect 21484 23780 21864 23832
rect 22058 23832 22192 23914
rect 22304 23862 22684 23914
rect 22304 23832 22438 23862
rect 22058 23780 22438 23832
rect 22550 23832 22684 23862
rect 22796 23862 23422 23914
rect 22796 23832 22930 23862
rect 22550 23780 22930 23832
rect 23042 23780 23176 23862
rect 23288 23780 23422 23862
rect 23616 23862 24242 23914
rect 23616 23780 23750 23862
rect 23862 23780 23996 23862
rect 24108 23832 24242 23862
rect 24354 23832 24488 23914
rect 24600 23832 24734 23914
rect 24846 23832 24980 23914
rect 24108 23780 24980 23832
rect 25174 23862 25554 23914
rect 25174 23780 25308 23862
rect 25420 23832 25554 23862
rect 25666 23862 26046 23914
rect 25666 23832 25800 23862
rect 25420 23780 25800 23832
rect 25912 23832 26046 23862
rect 26158 23832 26292 23914
rect 26404 23832 26538 23914
rect 26732 23832 26866 23914
rect 26978 23862 27850 23914
rect 26978 23832 27112 23862
rect 25912 23780 27112 23832
rect 27224 23780 27358 23862
rect 27470 23780 27604 23862
rect 27716 23832 27850 23862
rect 27962 23832 28178 23914
rect 28290 23862 28916 23914
rect 28290 23832 28424 23862
rect 27716 23780 28424 23832
rect 28536 23780 28670 23862
rect 28782 23832 28916 23862
rect 29028 23832 29162 23914
rect 29274 23862 30228 23914
rect 29274 23832 29408 23862
rect 28782 23780 29408 23832
rect 29602 23780 29736 23862
rect 29848 23780 29982 23862
rect 30094 23832 30228 23862
rect 30340 23832 30474 23914
rect 30586 23832 30720 23914
rect 30832 23832 30966 23914
rect 30094 23780 30966 23832
rect 31160 23832 31294 23914
rect 31406 23862 31786 23914
rect 31406 23832 31540 23862
rect 31160 23780 31540 23832
rect 31652 23780 31786 23862
rect 14268 23422 14402 23504
rect 31898 23422 32032 23504
rect 12710 23288 12844 23422
rect 13940 23370 14648 23422
rect 13940 23288 14074 23370
rect 14514 23340 14648 23370
rect 14760 23340 14894 23422
rect 15006 23370 15632 23422
rect 15006 23340 15140 23370
rect 14514 23288 15140 23340
rect 15252 23288 15386 23370
rect 15498 23340 15632 23370
rect 15744 23340 15878 23422
rect 16072 23370 18010 23422
rect 16072 23340 16206 23370
rect 15498 23288 16206 23340
rect 16318 23288 16452 23370
rect 16564 23288 16698 23370
rect 16810 23288 16944 23370
rect 17056 23288 17190 23370
rect 17302 23288 17518 23370
rect 17630 23288 17764 23370
rect 17876 23340 18010 23370
rect 18122 23340 18256 23422
rect 18368 23340 18502 23422
rect 18614 23370 19568 23422
rect 18614 23340 18748 23370
rect 17876 23288 18748 23340
rect 18942 23288 19076 23370
rect 19188 23288 19322 23370
rect 19434 23340 19568 23370
rect 19680 23370 20306 23422
rect 19680 23340 19814 23370
rect 19434 23288 19814 23340
rect 19926 23288 20060 23370
rect 20172 23340 20306 23370
rect 20500 23340 20634 23422
rect 20746 23370 21372 23422
rect 20746 23340 20880 23370
rect 20172 23288 20880 23340
rect 20992 23288 21126 23370
rect 21238 23340 21372 23370
rect 21484 23370 21864 23422
rect 21484 23340 21618 23370
rect 21238 23288 21618 23340
rect 21730 23340 21864 23370
rect 22058 23340 22192 23422
rect 22304 23370 22684 23422
rect 22304 23340 22438 23370
rect 21730 23288 22438 23340
rect 22550 23340 22684 23370
rect 22796 23340 22930 23422
rect 23042 23340 23176 23422
rect 23288 23370 23996 23422
rect 23288 23340 23422 23370
rect 22550 23288 23422 23340
rect 23616 23288 23750 23370
rect 23862 23340 23996 23370
rect 24108 23340 24242 23422
rect 24354 23370 25308 23422
rect 24354 23340 24488 23370
rect 23862 23288 24488 23340
rect 24600 23288 24734 23370
rect 24846 23288 24980 23370
rect 25174 23340 25308 23370
rect 25420 23370 26046 23422
rect 25420 23340 25554 23370
rect 25174 23288 25554 23340
rect 25666 23288 25800 23370
rect 25912 23340 26046 23370
rect 26158 23370 26538 23422
rect 26158 23340 26292 23370
rect 25912 23288 26292 23340
rect 26404 23340 26538 23370
rect 26732 23340 26866 23422
rect 26978 23340 27112 23422
rect 27224 23370 27604 23422
rect 27224 23340 27358 23370
rect 26404 23288 27358 23340
rect 27470 23340 27604 23370
rect 27716 23340 27850 23422
rect 27962 23340 28178 23422
rect 28290 23340 28424 23422
rect 28536 23340 28670 23422
rect 28782 23370 29162 23422
rect 28782 23340 28916 23370
rect 27470 23288 28916 23340
rect 29028 23340 29162 23370
rect 29274 23370 29982 23422
rect 29274 23340 29408 23370
rect 29028 23288 29408 23340
rect 29602 23288 29736 23370
rect 29848 23340 29982 23370
rect 30094 23370 30474 23422
rect 30094 23340 30228 23370
rect 29848 23288 30228 23340
rect 30340 23340 30474 23370
rect 30586 23370 30966 23422
rect 30586 23340 30720 23370
rect 30340 23288 30720 23340
rect 30832 23340 30966 23370
rect 31160 23340 31294 23422
rect 31406 23340 31540 23422
rect 31652 23370 32688 23422
rect 31652 23340 31786 23370
rect 30832 23288 31786 23340
rect 12710 22796 12844 22930
rect 13940 22878 14648 22930
rect 13940 22796 14074 22878
rect 14514 22796 14648 22878
rect 31652 22848 31786 22930
rect 31652 22796 32278 22848
rect 12710 22222 12844 22356
rect 13940 22274 14074 22356
rect 14514 22274 14648 22356
rect 13940 22222 14648 22274
rect 31652 22222 31786 22356
rect 12710 21730 12844 21864
rect 13940 21812 14648 21864
rect 13940 21730 14074 21812
rect 14514 21730 14648 21812
rect 31652 21812 32278 21864
rect 31652 21730 31786 21812
rect 12710 21238 12844 21372
rect 13940 21320 14648 21372
rect 13940 21290 14074 21320
rect 13858 21238 14074 21290
rect 14514 21238 14648 21320
rect 31652 21320 32688 21372
rect 31652 21238 31786 21320
rect 12710 20746 12844 20880
rect 13940 20798 14074 20880
rect 14514 20798 14648 20880
rect 13940 20746 14648 20798
rect 31652 20798 31786 20880
rect 31652 20746 32278 20798
rect 12710 20254 12844 20388
rect 13884 20336 14074 20388
rect 13940 20306 14074 20336
rect 14514 20306 14648 20388
rect 13940 20254 14648 20306
rect 31652 20306 31786 20388
rect 31652 20254 32688 20306
rect 12710 19680 12844 19814
rect 13940 19762 14648 19814
rect 13940 19680 14074 19762
rect 14514 19680 14648 19762
rect 31652 19762 32278 19814
rect 31652 19680 31786 19762
rect 12710 19188 12844 19322
rect 13940 19240 14074 19322
rect 14514 19240 14648 19322
rect 13940 19188 14648 19240
rect 31652 19240 31786 19322
rect 31652 19188 32688 19240
rect 12710 18696 12844 18830
rect 13940 18748 14074 18830
rect 14514 18748 14648 18830
rect 13940 18696 14648 18748
rect 31652 18748 31786 18830
rect 31652 18696 32278 18748
rect 12710 18204 12844 18338
rect 13940 18286 14648 18338
rect 13940 18256 14074 18286
rect 13940 18204 14156 18256
rect 14514 18204 14648 18286
rect 31652 18204 31786 18338
rect 12710 17712 12844 17846
rect 13940 17794 14648 17846
rect 13940 17712 14074 17794
rect 14514 17712 14648 17794
rect 31652 17794 32278 17846
rect 31652 17712 31786 17794
rect 12710 17190 12844 17272
rect 12628 17138 12844 17190
rect 13940 17220 14130 17272
rect 13940 17190 14074 17220
rect 14514 17190 14648 17272
rect 13940 17138 14648 17190
rect 31652 17190 31786 17272
rect 31652 17138 32688 17190
rect 12710 16646 12844 16780
rect 13940 16698 14074 16780
rect 14514 16698 14648 16780
rect 13940 16646 14648 16698
rect 31652 16728 32278 16780
rect 31652 16646 31786 16728
rect 8036 16154 8170 16288
rect 12654 16236 12844 16288
rect 12710 16206 12844 16236
rect 13940 16236 14648 16288
rect 12710 16154 12926 16206
rect 13940 16154 14074 16236
rect 14514 16154 14648 16236
rect 31652 16154 31786 16288
rect 7544 16042 7678 16124
rect 0 15990 7678 16042
rect 8508 16010 9169 16040
rect 8036 15796 8170 15878
rect 7980 15744 8170 15796
rect 12710 15662 12844 15796
rect 13940 15714 14074 15796
rect 14514 15714 14648 15796
rect 13940 15662 14648 15714
rect 31652 15714 31786 15796
rect 31652 15662 32278 15714
rect 7544 15550 7678 15632
rect 8508 15578 9103 15608
rect 0 15498 7678 15550
rect 8036 15334 8170 15468
rect 0 15252 7678 15304
rect 7544 15170 7678 15252
rect 12710 15252 12900 15304
rect 8508 15198 9037 15228
rect 12710 15170 12844 15252
rect 13940 15222 14074 15304
rect 14514 15222 14648 15304
rect 13940 15170 14648 15222
rect 31652 15170 31786 15304
rect 7954 15006 8170 15058
rect 8036 14924 8170 15006
rect 0 14760 7678 14812
rect 8508 14766 8971 14796
rect 7544 14678 7678 14760
rect 8036 14566 8170 14648
rect 12710 14596 12844 14730
rect 13940 14678 14648 14730
rect 13940 14596 14074 14678
rect 14514 14596 14648 14678
rect 31652 14678 32278 14730
rect 31652 14596 31786 14678
rect 8036 14514 9564 14566
rect 0 14432 7678 14484
rect 7593 14406 7645 14432
rect 8508 14386 8905 14416
rect 8750 14353 8816 14386
rect 8036 14186 9646 14238
rect 8036 14104 8170 14186
rect 9512 14156 9646 14186
rect 10332 14156 10466 14238
rect 9512 14104 10466 14156
rect 12710 14104 12844 14238
rect 13940 14186 14648 14238
rect 13940 14104 14074 14186
rect 14514 14104 14648 14186
rect 31652 14104 31786 14238
rect 9512 13664 9646 13746
rect 10332 13664 10466 13746
rect 9512 13612 10466 13664
rect 12710 13612 12844 13746
rect 13940 13664 14074 13746
rect 14514 13664 14648 13746
rect 13940 13612 14648 13664
rect 31652 13664 31786 13746
rect 31652 13612 32278 13664
rect 9512 13172 9646 13254
rect 10332 13172 10466 13254
rect 9512 13120 10466 13172
rect 12710 13172 12844 13254
rect 13940 13172 14074 13254
rect 14514 13172 14648 13254
rect 12710 13120 12926 13172
rect 13940 13120 14648 13172
rect 31652 13172 31786 13254
rect 31652 13120 32688 13172
rect 9512 12710 10466 12762
rect 9512 12628 9646 12710
rect 10332 12628 10466 12710
rect 12710 12680 12844 12762
rect 13940 12710 14648 12762
rect 13940 12680 14074 12710
rect 12710 12628 14074 12680
rect 14514 12628 14648 12710
rect 31652 12710 32278 12762
rect 31652 12628 31786 12710
rect 9512 12106 9646 12188
rect 10332 12106 10466 12188
rect 12710 12136 12900 12188
rect 12710 12106 12844 12136
rect 9512 12054 10466 12106
rect 12628 12054 12844 12106
rect 13940 12106 14074 12188
rect 14514 12106 14648 12188
rect 13940 12054 14648 12106
rect 31652 12054 31786 12188
rect 9512 11614 9646 11696
rect 10332 11614 10466 11696
rect 9512 11562 10466 11614
rect 12710 11562 12844 11696
rect 13940 11614 14074 11696
rect 14514 11614 14648 11696
rect 13940 11562 14648 11614
rect 31652 11614 31786 11696
rect 31652 11562 32278 11614
rect 9512 11152 10466 11204
rect 12654 11152 12844 11204
rect 9512 11070 9646 11152
rect 10332 11070 10466 11152
rect 12710 11070 12844 11152
rect 13940 11122 14074 11204
rect 14514 11122 14648 11204
rect 13940 11070 14648 11122
rect 31652 11122 31786 11204
rect 31652 11070 32688 11122
rect 9512 10660 10466 10712
rect 9512 10630 9646 10660
rect 9512 10578 9810 10630
rect 10332 10578 10466 10660
rect 12710 10578 12844 10712
rect 13940 10660 14648 10712
rect 13940 10578 14074 10660
rect 14514 10578 14648 10660
rect 31652 10660 32278 10712
rect 31652 10578 31786 10660
rect 9512 10138 9646 10220
rect 10332 10138 10466 10220
rect 12710 10138 12844 10220
rect 9512 10086 10466 10138
rect 12628 10086 12844 10138
rect 13940 10168 14648 10220
rect 13940 10086 14074 10168
rect 14514 10086 14648 10168
rect 31652 10086 31786 10220
rect 12710 9512 12844 9646
rect 13940 9564 14074 9646
rect 14514 9564 14648 9646
rect 13940 9512 14648 9564
rect 31652 9594 32278 9646
rect 31652 9512 31786 9594
rect 9758 9072 9892 9154
rect 10414 9072 10548 9154
rect 12654 9102 12844 9154
rect 12710 9072 12844 9102
rect 13940 9102 14648 9154
rect 13940 9072 14074 9102
rect 9758 9020 10548 9072
rect 12654 9020 12844 9072
rect 13884 9020 14074 9072
rect 14514 9020 14648 9102
rect 31652 9020 31786 9154
rect 9758 8580 9892 8662
rect 10414 8580 10548 8662
rect 9758 8528 10548 8580
rect 12710 8528 12844 8662
rect 13940 8580 14074 8662
rect 14514 8580 14648 8662
rect 13940 8528 14648 8580
rect 31652 8580 31786 8662
rect 31652 8528 32278 8580
rect 9758 8088 9892 8170
rect 10414 8088 10548 8170
rect 12628 8118 12844 8170
rect 13858 8118 14074 8170
rect 12710 8088 12844 8118
rect 1640 8006 1774 8088
rect 2296 8006 2430 8088
rect 9758 8036 10548 8088
rect 12628 8036 12844 8088
rect 13940 8088 14074 8118
rect 14514 8088 14648 8170
rect 13940 8036 14648 8088
rect 31652 8088 31786 8170
rect 31652 8036 32688 8088
rect 1640 7954 2430 8006
rect 1640 7596 1774 7678
rect 2296 7596 2430 7678
rect 1640 7544 2430 7596
rect 9758 7544 10548 7596
rect 9758 7514 9892 7544
rect 9758 7462 10384 7514
rect 10414 7462 10548 7544
rect 12710 7462 12844 7596
rect 13940 7544 14648 7596
rect 13940 7462 14074 7544
rect 14514 7462 14648 7544
rect 31652 7544 32278 7596
rect 31652 7462 31786 7544
rect 328 7216 1774 7268
rect 1640 7186 1774 7216
rect 2296 7186 2430 7268
rect 1640 7134 2512 7186
rect 9758 7052 10548 7104
rect 12654 7052 12844 7104
rect 9758 7022 9892 7052
rect 9758 6970 10302 7022
rect 10414 6970 10548 7052
rect 12710 6970 12844 7052
rect 13940 7052 14648 7104
rect 13940 7022 14074 7052
rect 13940 6970 14320 7022
rect 14514 6970 14648 7052
rect 31652 7022 31786 7104
rect 31514 6970 31786 7022
rect 1640 6806 2430 6858
rect 1640 6724 1774 6806
rect 2296 6724 2430 6806
rect 12792 6642 12926 6776
rect 12792 6612 12844 6642
rect 12710 6478 12844 6612
rect 14514 6560 14894 6612
rect 14514 6530 14648 6560
rect 14760 6530 14894 6560
rect 15006 6530 15140 6612
rect 15252 6530 15386 6612
rect 15498 6560 15878 6612
rect 15498 6530 15632 6560
rect 14514 6478 14730 6530
rect 14760 6478 15632 6530
rect 15744 6530 15878 6560
rect 16072 6560 16452 6612
rect 16072 6530 16206 6560
rect 15744 6478 16206 6530
rect 16318 6530 16452 6560
rect 16564 6530 16698 6612
rect 16810 6560 17190 6612
rect 16810 6530 16944 6560
rect 16318 6478 16944 6530
rect 17056 6530 17190 6560
rect 17302 6530 17518 6612
rect 17630 6530 17764 6612
rect 17876 6560 18502 6612
rect 17876 6530 18010 6560
rect 17056 6478 18010 6530
rect 18122 6478 18256 6560
rect 18368 6530 18502 6560
rect 18614 6530 18748 6612
rect 18942 6530 19076 6612
rect 19188 6530 19322 6612
rect 19434 6560 20060 6612
rect 19434 6530 19568 6560
rect 18368 6478 19568 6530
rect 19680 6478 19814 6560
rect 19926 6530 20060 6560
rect 20172 6560 20880 6612
rect 20172 6530 20306 6560
rect 19926 6478 20306 6530
rect 20500 6478 20634 6560
rect 20746 6530 20880 6560
rect 20992 6530 21126 6612
rect 21238 6530 21372 6612
rect 21484 6530 21618 6612
rect 21730 6560 22438 6612
rect 21730 6530 21864 6560
rect 20746 6478 21864 6530
rect 22058 6478 22192 6560
rect 22304 6530 22438 6560
rect 22550 6560 22930 6612
rect 22550 6530 22684 6560
rect 22304 6478 22684 6530
rect 22796 6530 22930 6560
rect 23042 6560 23422 6612
rect 23042 6530 23176 6560
rect 22796 6478 23176 6530
rect 23288 6530 23422 6560
rect 23616 6530 23750 6612
rect 23862 6530 23996 6612
rect 24108 6560 24734 6612
rect 24108 6530 24242 6560
rect 23288 6478 24242 6530
rect 24354 6478 24488 6560
rect 24600 6530 24734 6560
rect 24846 6530 24980 6612
rect 25174 6530 25308 6612
rect 25420 6530 25554 6612
rect 25666 6530 25800 6612
rect 25912 6560 26292 6612
rect 25912 6530 26046 6560
rect 24600 6478 26046 6530
rect 26158 6530 26292 6560
rect 26404 6530 26538 6612
rect 26732 6560 27358 6612
rect 26732 6530 26866 6560
rect 26158 6478 26866 6530
rect 26978 6478 27112 6560
rect 27224 6530 27358 6560
rect 27470 6560 29408 6612
rect 27470 6530 27604 6560
rect 27224 6478 27604 6530
rect 27716 6478 27850 6560
rect 27962 6478 28178 6560
rect 28290 6478 28424 6560
rect 28536 6478 28670 6560
rect 28782 6478 28916 6560
rect 29028 6478 29162 6560
rect 29274 6530 29408 6560
rect 29602 6530 29736 6612
rect 29848 6560 30228 6612
rect 29848 6530 29982 6560
rect 29274 6478 29982 6530
rect 30094 6530 30228 6560
rect 30340 6530 30474 6612
rect 30586 6530 30720 6612
rect 30832 6560 31540 6612
rect 30832 6530 30966 6560
rect 30094 6478 30966 6530
rect 31160 6478 31294 6560
rect 31406 6530 31540 6560
rect 31652 6530 31786 6612
rect 31406 6478 32278 6530
rect 1640 6366 1774 6448
rect 2296 6396 2486 6448
rect 2296 6366 2430 6396
rect 1640 6314 2430 6366
rect 14268 6120 14402 6202
rect 31898 6120 32032 6202
rect 14268 6068 14648 6120
rect 14514 6038 14648 6068
rect 14760 6038 14894 6120
rect 15006 6068 15386 6120
rect 15006 6038 15140 6068
rect 1640 5956 1774 6038
rect 2296 5956 2430 6038
rect 14514 5986 15140 6038
rect 15252 6038 15386 6068
rect 15498 6068 15878 6120
rect 15498 6038 15632 6068
rect 15252 5986 15632 6038
rect 15744 6038 15878 6068
rect 16072 6038 16206 6120
rect 16318 6038 16452 6120
rect 16564 6068 17190 6120
rect 16564 6038 16698 6068
rect 15744 5986 16698 6038
rect 16810 5986 16944 6068
rect 17056 6038 17190 6068
rect 17302 6068 18010 6120
rect 17302 6038 17518 6068
rect 17056 5986 17518 6038
rect 17630 5986 17764 6068
rect 17876 6038 18010 6068
rect 18122 6038 18256 6120
rect 18368 6068 18748 6120
rect 18368 6038 18502 6068
rect 17876 5986 18502 6038
rect 18614 6038 18748 6068
rect 18942 6038 19076 6120
rect 19188 6038 19322 6120
rect 19434 6068 19814 6120
rect 19434 6038 19568 6068
rect 18614 5986 19568 6038
rect 19680 6038 19814 6068
rect 19926 6068 20880 6120
rect 19926 6038 20060 6068
rect 19680 5986 20060 6038
rect 20172 5986 20306 6068
rect 20500 5986 20634 6068
rect 20746 6038 20880 6068
rect 20992 6038 21126 6120
rect 21238 6068 21864 6120
rect 21238 6038 21372 6068
rect 20746 5986 21372 6038
rect 21484 5986 21618 6068
rect 21730 6038 21864 6068
rect 22058 6038 22192 6120
rect 22304 6038 22438 6120
rect 22550 6038 22684 6120
rect 22796 6068 23422 6120
rect 22796 6038 22930 6068
rect 21730 5986 22930 6038
rect 23042 5986 23176 6068
rect 23288 6038 23422 6068
rect 23616 6068 24242 6120
rect 23616 6038 23750 6068
rect 23288 5986 23750 6038
rect 23862 5986 23996 6068
rect 24108 6038 24242 6068
rect 24354 6038 24488 6120
rect 24600 6038 24734 6120
rect 24846 6038 24980 6120
rect 25174 6068 25554 6120
rect 25174 6038 25308 6068
rect 24108 5986 25308 6038
rect 25420 6038 25554 6068
rect 25666 6038 25800 6120
rect 25912 6038 26046 6120
rect 26158 6068 26538 6120
rect 26158 6038 26292 6068
rect 25420 5986 26292 6038
rect 26404 6038 26538 6068
rect 26732 6038 26866 6120
rect 26978 6068 27850 6120
rect 26978 6038 27112 6068
rect 26404 5986 27112 6038
rect 27224 5986 27358 6068
rect 27470 5986 27604 6068
rect 27716 6038 27850 6068
rect 27962 6038 28178 6120
rect 28290 6038 28424 6120
rect 28536 6068 28916 6120
rect 28536 6038 28670 6068
rect 27716 5986 28670 6038
rect 28782 6038 28916 6068
rect 29028 6068 29736 6120
rect 29028 6038 29162 6068
rect 28782 5986 29162 6038
rect 29274 5986 29408 6068
rect 29602 6038 29736 6068
rect 29848 6068 30228 6120
rect 29848 6038 29982 6068
rect 29602 5986 29982 6038
rect 30094 6038 30228 6068
rect 30340 6038 30474 6120
rect 30586 6038 30720 6120
rect 30832 6038 30966 6120
rect 31160 6038 31294 6120
rect 31406 6068 32688 6120
rect 31406 6038 31540 6068
rect 30094 5986 31540 6038
rect 31652 5986 31786 6068
rect 1640 5904 2430 5956
rect 14704 5822 14976 5874
rect 14842 5792 14976 5822
rect 15088 5792 15222 5874
rect 15334 5792 15468 5874
rect 15580 5822 15960 5874
rect 15580 5792 15714 5822
rect 8750 5756 12945 5786
rect 14842 5740 15714 5792
rect 15826 5792 15960 5822
rect 16154 5792 16288 5874
rect 16400 5822 16780 5874
rect 16400 5792 16534 5822
rect 15826 5740 16534 5792
rect 16646 5792 16780 5822
rect 16892 5792 17026 5874
rect 17138 5792 17272 5874
rect 17384 5792 17518 5874
rect 17712 5792 17846 5874
rect 17958 5822 18338 5874
rect 17958 5792 18092 5822
rect 16646 5740 18092 5792
rect 18204 5792 18338 5822
rect 18450 5822 18830 5874
rect 18450 5792 18584 5822
rect 18204 5740 18584 5792
rect 18696 5792 18830 5822
rect 18942 5792 19158 5874
rect 19270 5822 19650 5874
rect 19270 5792 19404 5822
rect 18696 5740 19404 5792
rect 19516 5792 19650 5822
rect 19762 5792 19896 5874
rect 20008 5822 20716 5874
rect 20008 5792 20142 5822
rect 19516 5740 20142 5792
rect 20254 5740 20388 5822
rect 20582 5792 20716 5822
rect 20828 5792 20962 5874
rect 21074 5792 21208 5874
rect 21320 5792 21454 5874
rect 21566 5792 21700 5874
rect 21812 5822 22274 5874
rect 21812 5792 21946 5822
rect 20582 5740 21946 5792
rect 22140 5792 22274 5822
rect 22386 5822 23258 5874
rect 22386 5792 22520 5822
rect 22140 5740 22520 5792
rect 22632 5740 22766 5822
rect 22878 5740 23012 5822
rect 23124 5792 23258 5822
rect 23370 5792 23504 5874
rect 23698 5822 24078 5874
rect 23698 5792 23832 5822
rect 23124 5740 23832 5792
rect 23944 5792 24078 5822
rect 24190 5822 25062 5874
rect 24190 5792 24324 5822
rect 23944 5740 24324 5792
rect 24436 5740 24570 5822
rect 24682 5740 24816 5822
rect 24928 5792 25062 5822
rect 25256 5792 25390 5874
rect 25502 5792 25636 5874
rect 25748 5792 25882 5874
rect 25994 5792 26128 5874
rect 26240 5822 26620 5874
rect 26240 5792 26374 5822
rect 24928 5740 26374 5792
rect 26486 5792 26620 5822
rect 26814 5792 26948 5874
rect 27060 5822 27440 5874
rect 27060 5792 27194 5822
rect 26486 5740 27194 5792
rect 27306 5792 27440 5822
rect 27552 5792 27686 5874
rect 27798 5792 27932 5874
rect 28044 5792 28178 5874
rect 28372 5792 28506 5874
rect 28618 5822 28998 5874
rect 28618 5792 28752 5822
rect 27306 5740 28752 5792
rect 28864 5792 28998 5822
rect 29110 5822 29490 5874
rect 29110 5792 29244 5822
rect 28864 5740 29244 5792
rect 29356 5792 29490 5822
rect 29602 5792 29818 5874
rect 29930 5792 30064 5874
rect 30176 5792 30310 5874
rect 30422 5792 30556 5874
rect 30668 5822 31376 5874
rect 30668 5792 30802 5822
rect 29356 5740 30802 5792
rect 30914 5740 31048 5822
rect 31242 5792 31376 5822
rect 31488 5792 31622 5874
rect 31242 5740 31622 5792
rect 1640 5576 2430 5628
rect 10276 5576 10466 5628
rect 1640 5546 1774 5576
rect 1640 5494 1856 5546
rect 2296 5494 2430 5576
rect 10332 5546 10466 5576
rect 10276 5494 10466 5546
rect 11316 5494 11450 5628
rect 1640 5166 2430 5218
rect 10332 5166 10466 5218
rect 11316 5166 11450 5218
rect 1688 5121 1740 5166
rect 2316 5121 2368 5166
rect 10362 5101 10414 5166
rect 11332 5101 11384 5166
rect 1201 5046 14746 5076
rect 8750 4943 13927 4973
rect 1640 4756 1830 4808
rect 1640 4726 1774 4756
rect 2296 4726 2430 4808
rect 10250 4756 10466 4808
rect 1640 4674 2430 4726
rect 10332 4674 10466 4756
rect 11316 4674 11450 4808
rect 15170 4562 15304 4644
rect 15416 4562 15550 4644
rect 15662 4562 15796 4644
rect 15908 4592 16288 4644
rect 15908 4562 16042 4592
rect 8750 4508 14091 4538
rect 15170 4510 16042 4562
rect 16154 4562 16288 4592
rect 16400 4562 16534 4644
rect 16728 4592 17354 4644
rect 16728 4562 16862 4592
rect 16154 4510 16862 4562
rect 16974 4510 17108 4592
rect 17220 4562 17354 4592
rect 17466 4592 17846 4644
rect 17466 4562 17600 4592
rect 17220 4510 17600 4562
rect 17712 4562 17846 4592
rect 17958 4562 18092 4644
rect 18286 4592 18666 4644
rect 18286 4562 18420 4592
rect 17712 4510 18420 4562
rect 18532 4562 18666 4592
rect 18778 4562 18912 4644
rect 19024 4562 19158 4644
rect 19270 4562 19404 4644
rect 19516 4592 19978 4644
rect 19516 4562 19650 4592
rect 18532 4510 19650 4562
rect 19844 4562 19978 4592
rect 20090 4592 20470 4644
rect 20090 4562 20224 4592
rect 19844 4510 20224 4562
rect 20336 4562 20470 4592
rect 20582 4592 20962 4644
rect 20582 4562 20716 4592
rect 20336 4510 20716 4562
rect 20828 4562 20962 4592
rect 21074 4592 21536 4644
rect 21074 4562 21208 4592
rect 20828 4510 21208 4562
rect 21402 4562 21536 4592
rect 21648 4592 22028 4644
rect 21648 4562 21782 4592
rect 21402 4510 21782 4562
rect 21894 4562 22028 4592
rect 22140 4592 22520 4644
rect 22140 4562 22274 4592
rect 21894 4510 22274 4562
rect 22386 4562 22520 4592
rect 22632 4562 22848 4644
rect 22960 4592 23586 4644
rect 22960 4562 23094 4592
rect 22386 4510 23094 4562
rect 23206 4510 23340 4592
rect 23452 4562 23586 4592
rect 23698 4562 23832 4644
rect 23944 4562 24078 4644
rect 24272 4562 24406 4644
rect 24518 4592 24898 4644
rect 24518 4562 24652 4592
rect 23452 4510 24652 4562
rect 24764 4562 24898 4592
rect 25010 4592 25390 4644
rect 25010 4562 25144 4592
rect 24764 4510 25144 4562
rect 25256 4562 25390 4592
rect 25502 4592 25964 4644
rect 25502 4562 25636 4592
rect 25256 4510 25636 4562
rect 25830 4562 25964 4592
rect 26076 4562 26210 4644
rect 26322 4562 26456 4644
rect 26568 4592 26948 4644
rect 26568 4562 26702 4592
rect 25830 4510 26702 4562
rect 26814 4562 26948 4592
rect 27060 4562 27194 4644
rect 27388 4592 27768 4644
rect 27388 4562 27522 4592
rect 26814 4510 27522 4562
rect 27634 4562 27768 4592
rect 27880 4592 28260 4644
rect 27880 4562 28014 4592
rect 27634 4510 28014 4562
rect 28126 4562 28260 4592
rect 28372 4592 28752 4644
rect 28372 4562 28506 4592
rect 28126 4510 28506 4562
rect 28618 4562 28752 4592
rect 28946 4592 29572 4644
rect 28946 4562 29080 4592
rect 28618 4510 29080 4562
rect 29192 4510 29326 4592
rect 29438 4562 29572 4592
rect 29684 4562 29818 4644
rect 29930 4592 30638 4644
rect 29930 4562 30064 4592
rect 29438 4510 30064 4562
rect 30176 4510 30310 4592
rect 30504 4562 30638 4592
rect 30750 4592 31130 4644
rect 30750 4562 30884 4592
rect 30504 4510 30884 4562
rect 30996 4562 31130 4592
rect 31242 4592 31622 4644
rect 31242 4562 31376 4592
rect 30996 4510 31376 4562
rect 31488 4562 31622 4592
rect 31488 4510 32688 4562
rect 1640 4346 2430 4398
rect 1640 4316 1774 4346
rect 738 4264 1774 4316
rect 2296 4264 2430 4346
rect 10332 4264 10466 4398
rect 11316 4264 11450 4398
rect 8750 4131 14009 4161
rect 10332 3906 10466 3988
rect 10332 3854 10522 3906
rect 11316 3854 11450 3988
rect 984 3496 1118 3578
rect 328 3444 1118 3496
rect 10332 3444 10466 3578
rect 11316 3444 11450 3578
rect 0 3280 1282 3332
rect 1148 3198 1282 3280
rect 15170 3250 15304 3332
rect 17220 3250 17354 3332
rect 19270 3250 19404 3332
rect 21402 3250 21536 3332
rect 23452 3250 23586 3332
rect 25584 3250 25718 3332
rect 27634 3250 27768 3332
rect 29684 3250 29818 3332
rect 15170 3198 15714 3250
rect 17220 3198 17764 3250
rect 19270 3198 19814 3250
rect 21402 3198 21946 3250
rect 23452 3198 23996 3250
rect 25584 3198 26046 3250
rect 27634 3198 28096 3250
rect 29684 3198 30228 3250
rect 984 3086 1118 3168
rect 10332 3116 10548 3168
rect 10332 3086 10466 3116
rect 738 3034 1118 3086
rect 10276 3034 10466 3086
rect 11316 3034 11450 3168
rect 15416 3004 15550 3086
rect 1148 2922 1282 3004
rect 0 2870 1282 2922
rect 4182 2870 4316 3004
rect 15416 2952 15632 3004
rect 17466 2952 17600 3086
rect 19598 2952 19732 3086
rect 21648 2952 21782 3086
rect 23698 2952 23832 3086
rect 25830 2952 25964 3086
rect 27880 2952 28014 3086
rect 30012 3004 30146 3086
rect 30012 2952 33016 3004
rect 15170 2758 15304 2840
rect 17220 2758 17354 2840
rect 19270 2758 19404 2840
rect 21402 2758 21536 2840
rect 23452 2758 23586 2840
rect 25584 2758 25718 2840
rect 27634 2758 27768 2840
rect 29684 2758 29818 2840
rect 984 2624 1118 2758
rect 10332 2676 10466 2758
rect 11316 2676 11450 2758
rect 15170 2706 15550 2758
rect 17220 2706 17846 2758
rect 19270 2706 19896 2758
rect 21402 2706 21618 2758
rect 23452 2706 24078 2758
rect 25584 2706 26128 2758
rect 27634 2706 28178 2758
rect 29684 2706 30310 2758
rect 10332 2624 11450 2676
rect 15580 2594 15714 2676
rect 15580 2542 16288 2594
rect 17712 2542 17846 2676
rect 19762 2542 19896 2676
rect 21812 2624 23504 2676
rect 23944 2624 25636 2676
rect 25994 2624 27686 2676
rect 28044 2624 29736 2676
rect 21812 2594 21946 2624
rect 21812 2542 22110 2594
rect 23944 2542 24078 2624
rect 25994 2542 26128 2624
rect 28044 2542 28178 2624
rect 30176 2542 30310 2676
rect 10250 2296 11450 2348
rect 10332 2266 10466 2296
rect 10332 2214 10548 2266
rect 11316 2214 11450 2296
rect 15524 2050 15714 2102
rect 15580 1968 15714 2050
rect 17712 2020 17846 2102
rect 17656 1968 17846 2020
rect 19762 1968 19896 2102
rect 21592 2050 23586 2102
rect 21812 2020 21946 2050
rect 21812 1968 22028 2020
rect 23944 1968 24078 2102
rect 25994 1968 26128 2102
rect 28044 2050 29818 2102
rect 28044 1968 28178 2050
rect 30176 1968 30310 2102
rect 10414 1476 10548 1528
rect 10414 1364 10471 1476
rect 9922 1312 10056 1364
rect 10414 1312 10548 1364
rect 11070 1312 11204 1364
rect 11562 1312 11696 1528
rect 12218 1312 12352 1364
rect 12710 1312 12844 1528
rect 13366 1312 13500 1364
rect 13858 1312 13992 1528
rect 15006 1476 15140 1528
rect 15078 1364 15140 1476
rect 16236 1476 16370 1528
rect 17384 1476 17764 1528
rect 16236 1364 16296 1476
rect 17384 1364 17518 1476
rect 14514 1312 14648 1364
rect 15006 1312 15140 1364
rect 15744 1312 15878 1364
rect 16236 1312 16370 1364
rect 16892 1312 17026 1364
rect 17302 1312 17518 1364
rect 18040 1312 18174 1364
rect 18532 1312 18666 1528
rect 19188 1312 19322 1364
rect 19680 1312 19814 1528
rect 20828 1476 20962 1528
rect 20904 1364 20962 1476
rect 22058 1476 22192 1528
rect 22058 1364 22120 1476
rect 20336 1312 20470 1364
rect 20828 1312 20962 1364
rect 21566 1312 21700 1364
rect 22058 1312 22192 1364
rect 9923 1235 9975 1312
rect 11088 1235 11140 1312
rect 12253 1235 12305 1312
rect 13418 1235 13470 1312
rect 14583 1235 14635 1312
rect 15748 1235 15800 1312
rect 16913 1235 16965 1312
rect 18078 1235 18130 1312
rect 19243 1235 19295 1312
rect 20408 1235 20460 1312
rect 21573 1235 21625 1312
rect 8816 1193 11662 1223
rect 10414 984 10548 1118
rect 11562 984 11696 1118
rect 12710 984 12844 1118
rect 13858 984 13992 1118
rect 15006 1066 15714 1118
rect 15006 984 15140 1066
rect 16236 984 16370 1118
rect 17384 1066 17682 1118
rect 17384 1036 17518 1066
rect 17384 984 17682 1036
rect 18532 984 18666 1118
rect 19680 1066 19896 1118
rect 19680 1036 19814 1066
rect 19598 984 19814 1036
rect 20828 984 20962 1118
rect 22002 1066 22192 1118
rect 22058 984 22192 1066
rect 574 574 32442 790
rect 164 164 32852 380
<< metal4 >>
rect 164 164 380 24734
rect 574 574 790 24324
rect 12710 23396 12762 24570
rect 14514 23888 14566 24160
rect 16072 23888 16124 24160
rect 20500 23888 20552 24160
rect 22878 23888 22930 24160
rect 23944 23888 23996 24160
rect 25174 23888 25226 24160
rect 31160 23888 31212 24160
rect 12710 21812 12762 22822
rect 12792 22304 12844 23314
rect 14022 22904 14074 23832
rect 14514 22330 14566 23340
rect 12710 20854 12762 21782
rect 12792 21320 12844 22248
rect 12710 19762 12762 20772
rect 12792 20362 12844 21290
rect 13858 20336 13910 21264
rect 13940 20854 13992 21782
rect 14022 21346 14074 22274
rect 31734 21346 31786 22274
rect 12710 18778 12762 19706
rect 12792 19296 12844 20306
rect 13940 19270 13992 20280
rect 14022 19762 14074 20772
rect 12710 17820 12762 18748
rect 12792 18286 12844 19214
rect 12628 16236 12680 17164
rect 12710 16728 12762 17738
rect 12792 17246 12844 18256
rect 14022 17794 14074 18722
rect 14514 18286 14566 19214
rect 14596 18804 14648 19732
rect 31734 18286 31786 19214
rect 13940 16728 13992 17738
rect 14104 17220 14156 18230
rect 7954 15032 8006 15796
rect 8118 15416 8170 16180
rect 12792 15770 12844 16698
rect 8036 14596 8088 15360
rect 8118 14186 8170 14950
rect 12710 14678 12762 15688
rect 12874 15252 12926 16180
rect 13940 15770 13992 16698
rect 14022 16262 14074 17190
rect 31734 16236 31786 17164
rect 14022 15278 14074 16206
rect 9512 13694 9564 14540
rect 9594 13228 9646 14156
rect 12710 13694 12762 14622
rect 12792 14212 12844 15222
rect 10332 12736 10384 13664
rect 9512 11152 9564 12080
rect 9594 11670 9646 12680
rect 10414 12136 10466 13146
rect 12710 12736 12762 13664
rect 12792 13202 12844 14130
rect 13940 13720 13992 14648
rect 14022 14212 14074 15222
rect 14596 14678 14648 15688
rect 31734 15252 31786 16180
rect 9512 10194 9564 11122
rect 9594 10660 9646 11588
rect 12628 11152 12680 12080
rect 12792 11644 12844 12654
rect 12874 12136 12926 13146
rect 13940 11644 13992 12654
rect 14022 12162 14074 13172
rect 14514 12736 14566 13664
rect 14596 13202 14648 14130
rect 31652 13202 31704 14130
rect 12710 10660 12762 11588
rect 9758 8610 9810 10604
rect 10414 9102 10466 10112
rect 12628 9102 12680 10112
rect 12710 9620 12762 10630
rect 12792 10194 12844 11122
rect 13940 10686 13992 11614
rect 14514 11152 14566 12080
rect 31734 11178 31786 12106
rect 13940 9594 13992 10604
rect 14022 10194 14074 11122
rect 31734 10168 31786 11096
rect 1186 5061 1216 7797
rect 1640 7242 1692 8006
rect 2296 6832 2348 7596
rect 9758 7544 9810 8554
rect 9840 8118 9892 9046
rect 12628 8144 12680 9072
rect 12792 8610 12844 9538
rect 1640 5192 1692 5956
rect 1722 5602 1774 6366
rect 2378 6012 2430 6776
rect 2460 6396 2512 7160
rect 9840 7052 9892 8062
rect 10250 5576 10302 6996
rect 1722 4372 1774 5218
rect 1804 4756 1856 5520
rect 10250 4782 10302 5546
rect 10332 5166 10384 7488
rect 12628 7052 12680 8062
rect 12710 7544 12762 8554
rect 13858 8144 13910 9072
rect 13940 8636 13992 9564
rect 12792 6724 12844 7488
rect 13940 7078 13992 8088
rect 14022 7544 14074 8554
rect 31652 8118 31704 9046
rect 14268 6150 14320 6996
rect 14596 6560 14648 7488
rect 14678 5822 14730 6504
rect 31488 6094 31540 7022
rect 10332 3936 10384 4700
rect 10414 4346 10466 5192
rect 11316 4346 11368 5192
rect 11398 4782 11450 5546
rect 10414 3552 10466 4316
rect 1066 2732 1118 3496
rect 4182 0 4234 2896
rect 10250 2322 10302 3086
rect 10332 2732 10384 3496
rect 10496 3142 10548 3906
rect 11316 3552 11368 4316
rect 11398 3962 11450 4726
rect 11316 2732 11368 3496
rect 11398 3116 11450 3880
rect 10414 1476 10466 2650
rect 11398 2322 11450 3086
rect 9922 0 9974 1338
rect 10414 738 10466 1338
rect 10496 1066 10548 2240
rect 15498 2050 15550 2732
rect 10496 328 10548 1010
rect 11152 0 11204 1338
rect 11562 738 11614 1338
rect 11644 328 11696 1010
rect 12300 0 12352 1338
rect 12710 738 12762 1338
rect 12792 328 12844 1010
rect 13448 0 13500 1338
rect 13858 738 13910 1338
rect 13940 328 13992 1010
rect 14596 0 14648 1338
rect 15006 738 15058 1338
rect 15088 328 15140 1010
rect 15580 0 15632 2978
rect 15662 2624 15714 3224
rect 15662 1092 15714 2020
rect 16236 1476 16288 2568
rect 15744 0 15796 1338
rect 16236 738 16288 1338
rect 16318 328 16370 1010
rect 16974 0 17026 1338
rect 17302 738 17354 1338
rect 17466 0 17518 2978
rect 17712 2624 17764 3224
rect 17630 1092 17682 2020
rect 17712 1502 17764 2594
rect 17794 2050 17846 2732
rect 17630 328 17682 1010
rect 18040 0 18092 1338
rect 18532 738 18584 1338
rect 18614 328 18666 1010
rect 19270 0 19322 1338
rect 19598 328 19650 1010
rect 19680 0 19732 2978
rect 19762 2624 19814 3224
rect 19762 1502 19814 2594
rect 19844 2050 19896 2732
rect 21566 2050 21618 2732
rect 19762 738 19814 1338
rect 19844 1092 19896 2020
rect 20418 0 20470 1338
rect 20828 328 20880 1010
rect 20910 738 20962 1338
rect 21566 0 21618 1338
rect 21730 0 21782 2978
rect 21894 2624 21946 3224
rect 23452 2650 23504 3250
rect 21976 1066 22028 1994
rect 22058 1476 22110 2568
rect 23534 2076 23586 2758
rect 22058 328 22110 1010
rect 22140 738 22192 1338
rect 23780 0 23832 2978
rect 23944 2624 23996 3224
rect 24026 2050 24078 2732
rect 25584 2650 25636 3250
rect 25912 0 25964 2978
rect 25994 2624 26046 3224
rect 26076 2050 26128 2732
rect 27634 2650 27686 3250
rect 25994 328 26046 1994
rect 27880 0 27932 2978
rect 28044 2624 28096 3224
rect 28126 2050 28178 2732
rect 29684 2650 29736 3250
rect 29766 2076 29818 2758
rect 30176 2624 30228 3224
rect 30258 2050 30310 2732
rect 28126 328 28178 1994
rect 32226 574 32442 24324
rect 32636 164 32852 24734
use bank  bank_0
timestamp 1574592810
transform 1 0 8882 0 1 1912
box 0 0 23074 21989
use col_addr_dff  col_addr_dff_0
timestamp 1574592812
transform 1 0 9915 0 1 1014
box -116 -36 3495 451
use contact_6  contact_6_0
timestamp 1574592811
transform 1 0 30016 0 1 3018
box 0 0 46 46
use contact_6  contact_6_1
timestamp 1574592811
transform 1 0 27936 0 1 3018
box 0 0 46 46
use contact_6  contact_6_2
timestamp 1574592811
transform 1 0 25856 0 1 3018
box 0 0 46 46
use contact_6  contact_6_3
timestamp 1574592811
transform 1 0 23776 0 1 3018
box 0 0 46 46
use contact_6  contact_6_4
timestamp 1574592811
transform 1 0 21696 0 1 3018
box 0 0 46 46
use contact_6  contact_6_5
timestamp 1574592811
transform 1 0 19616 0 1 3018
box 0 0 46 46
use contact_6  contact_6_6
timestamp 1574592811
transform 1 0 17536 0 1 3018
box 0 0 46 46
use contact_6  contact_6_7
timestamp 1574592811
transform 1 0 15456 0 1 3018
box 0 0 46 46
use contact_7  contact_7_0
timestamp 1574592811
transform 1 0 7593 0 1 16030
box 0 0 52 52
use contact_7  contact_7_1
timestamp 1574592811
transform 1 0 7593 0 1 15536
box 0 0 52 52
use contact_7  contact_7_2
timestamp 1574592811
transform 1 0 7593 0 1 15218
box 0 0 52 52
use contact_7  contact_7_3
timestamp 1574592811
transform 1 0 7593 0 1 14724
box 0 0 52 52
use contact_7  contact_7_4
timestamp 1574592811
transform 1 0 7593 0 1 14406
box 0 0 52 52
use contact_7  contact_7_5
timestamp 1574592811
transform 1 0 12253 0 1 1235
box 0 0 52 52
use contact_7  contact_7_6
timestamp 1574592811
transform 1 0 11088 0 1 1235
box 0 0 52 52
use contact_7  contact_7_7
timestamp 1574592811
transform 1 0 9923 0 1 1235
box 0 0 52 52
use contact_7  contact_7_8
timestamp 1574592811
transform 1 0 30013 0 1 3016
box 0 0 52 52
use contact_7  contact_7_9
timestamp 1574592811
transform 1 0 27933 0 1 3016
box 0 0 52 52
use contact_7  contact_7_10
timestamp 1574592811
transform 1 0 25853 0 1 3016
box 0 0 52 52
use contact_7  contact_7_11
timestamp 1574592811
transform 1 0 23773 0 1 3016
box 0 0 52 52
use contact_7  contact_7_12
timestamp 1574592811
transform 1 0 21693 0 1 3016
box 0 0 52 52
use contact_7  contact_7_13
timestamp 1574592811
transform 1 0 19613 0 1 3016
box 0 0 52 52
use contact_7  contact_7_14
timestamp 1574592811
transform 1 0 17533 0 1 3016
box 0 0 52 52
use contact_7  contact_7_15
timestamp 1574592811
transform 1 0 15453 0 1 3016
box 0 0 52 52
use contact_7  contact_7_16
timestamp 1574592811
transform 1 0 21573 0 1 1235
box 0 0 52 52
use contact_7  contact_7_17
timestamp 1574592811
transform 1 0 20408 0 1 1235
box 0 0 52 52
use contact_7  contact_7_18
timestamp 1574592811
transform 1 0 19243 0 1 1235
box 0 0 52 52
use contact_7  contact_7_19
timestamp 1574592811
transform 1 0 18078 0 1 1235
box 0 0 52 52
use contact_7  contact_7_20
timestamp 1574592811
transform 1 0 16913 0 1 1235
box 0 0 52 52
use contact_7  contact_7_21
timestamp 1574592811
transform 1 0 15748 0 1 1235
box 0 0 52 52
use contact_7  contact_7_22
timestamp 1574592811
transform 1 0 14583 0 1 1235
box 0 0 52 52
use contact_7  contact_7_23
timestamp 1574592811
transform 1 0 13418 0 1 1235
box 0 0 52 52
use contact_7  contact_7_24
timestamp 1574592811
transform 1 0 4259 0 1 2877
box 0 0 52 52
use contact_7  contact_7_25
timestamp 1574592811
transform 1 0 1154 0 1 3250
box 0 0 52 52
use contact_7  contact_7_26
timestamp 1574592811
transform 1 0 1154 0 1 2932
box 0 0 52 52
use contact_7  contact_7_27
timestamp 1574592811
transform 1 0 9143 0 1 15999
box 0 0 52 52
use contact_7  contact_7_28
timestamp 1574592811
transform 1 0 8482 0 1 15999
box 0 0 52 52
use contact_7  contact_7_29
timestamp 1574592811
transform 1 0 9077 0 1 15567
box 0 0 52 52
use contact_7  contact_7_30
timestamp 1574592811
transform 1 0 8482 0 1 15567
box 0 0 52 52
use contact_7  contact_7_31
timestamp 1574592811
transform 1 0 9011 0 1 15187
box 0 0 52 52
use contact_7  contact_7_32
timestamp 1574592811
transform 1 0 8482 0 1 15187
box 0 0 52 52
use contact_7  contact_7_33
timestamp 1574592811
transform 1 0 8945 0 1 14755
box 0 0 52 52
use contact_7  contact_7_34
timestamp 1574592811
transform 1 0 8482 0 1 14755
box 0 0 52 52
use contact_7  contact_7_35
timestamp 1574592811
transform 1 0 8879 0 1 14375
box 0 0 52 52
use contact_7  contact_7_36
timestamp 1574592811
transform 1 0 8482 0 1 14375
box 0 0 52 52
use contact_7  contact_7_37
timestamp 1574592811
transform 1 0 1175 0 1 7771
box 0 0 52 52
use contact_7  contact_7_38
timestamp 1574592811
transform 1 0 12919 0 1 5745
box 0 0 52 52
use contact_7  contact_7_39
timestamp 1574592811
transform 1 0 8724 0 1 5745
box 0 0 52 52
use contact_7  contact_7_40
timestamp 1574592811
transform 1 0 13901 0 1 4932
box 0 0 52 52
use contact_7  contact_7_41
timestamp 1574592811
transform 1 0 8724 0 1 4932
box 0 0 52 52
use contact_7  contact_7_42
timestamp 1574592811
transform 1 0 14065 0 1 4497
box 0 0 52 52
use contact_7  contact_7_43
timestamp 1574592811
transform 1 0 8724 0 1 4497
box 0 0 52 52
use contact_7  contact_7_44
timestamp 1574592811
transform 1 0 13983 0 1 4120
box 0 0 52 52
use contact_7  contact_7_45
timestamp 1574592811
transform 1 0 8724 0 1 4120
box 0 0 52 52
use contact_16  contact_16_0
timestamp 1574592811
transform 1 0 30024 0 1 3027
box 0 0 29 29
use contact_16  contact_16_1
timestamp 1574592811
transform 1 0 27944 0 1 3027
box 0 0 29 29
use contact_16  contact_16_2
timestamp 1574592811
transform 1 0 25864 0 1 3027
box 0 0 29 29
use contact_16  contact_16_3
timestamp 1574592811
transform 1 0 23784 0 1 3027
box 0 0 29 29
use contact_16  contact_16_4
timestamp 1574592811
transform 1 0 21704 0 1 3027
box 0 0 29 29
use contact_16  contact_16_5
timestamp 1574592811
transform 1 0 19624 0 1 3027
box 0 0 29 29
use contact_16  contact_16_6
timestamp 1574592811
transform 1 0 17544 0 1 3027
box 0 0 29 29
use contact_16  contact_16_7
timestamp 1574592811
transform 1 0 15464 0 1 3027
box 0 0 29 29
use contact_30  contact_30_0
timestamp 1574592812
transform 1 0 8790 0 1 1182
box 0 0 52 52
use contact_30  contact_30_1
timestamp 1574592812
transform 1 0 8790 0 1 14353
box 0 0 52 52
use contact_32  contact_32_0
timestamp 1574592813
transform 1 0 32636 0 1 6068
box 0 0 52 52
use contact_32  contact_32_1
timestamp 1574592813
transform 1 0 32636 0 1 23370
box 0 0 52 52
use contact_32  contact_32_2
timestamp 1574592813
transform 1 0 32636 0 1 13120
box 0 0 52 52
use contact_32  contact_32_3
timestamp 1574592813
transform 1 0 31652 0 1 13202
box 0 0 52 52
use contact_32  contact_32_4
timestamp 1574592813
transform 1 0 31652 0 1 14104
box 0 0 52 52
use contact_32  contact_32_5
timestamp 1574592813
transform 1 0 32636 0 1 8036
box 0 0 52 52
use contact_32  contact_32_6
timestamp 1574592813
transform 1 0 32636 0 1 19188
box 0 0 52 52
use contact_32  contact_32_7
timestamp 1574592813
transform 1 0 31734 0 1 18286
box 0 0 52 52
use contact_32  contact_32_8
timestamp 1574592813
transform 1 0 31734 0 1 19188
box 0 0 52 52
use contact_32  contact_32_9
timestamp 1574592813
transform 1 0 31652 0 1 8118
box 0 0 52 52
use contact_32  contact_32_10
timestamp 1574592813
transform 1 0 31652 0 1 9020
box 0 0 52 52
use contact_32  contact_32_11
timestamp 1574592813
transform 1 0 32636 0 1 20254
box 0 0 52 52
use contact_32  contact_32_12
timestamp 1574592813
transform 1 0 31734 0 1 15252
box 0 0 52 52
use contact_32  contact_32_13
timestamp 1574592813
transform 1 0 31734 0 1 16154
box 0 0 52 52
use contact_32  contact_32_14
timestamp 1574592813
transform 1 0 32636 0 1 21320
box 0 0 52 52
use contact_32  contact_32_15
timestamp 1574592813
transform 1 0 31734 0 1 22222
box 0 0 52 52
use contact_32  contact_32_16
timestamp 1574592813
transform 1 0 31734 0 1 21320
box 0 0 52 52
use contact_32  contact_32_17
timestamp 1574592813
transform 1 0 32636 0 1 11070
box 0 0 52 52
use contact_32  contact_32_18
timestamp 1574592813
transform 1 0 31734 0 1 10168
box 0 0 52 52
use contact_32  contact_32_19
timestamp 1574592813
transform 1 0 31734 0 1 11070
box 0 0 52 52
use contact_32  contact_32_20
timestamp 1574592813
transform 1 0 31734 0 1 12054
box 0 0 52 52
use contact_32  contact_32_21
timestamp 1574592813
transform 1 0 31734 0 1 11152
box 0 0 52 52
use contact_32  contact_32_22
timestamp 1574592813
transform 1 0 32636 0 1 17138
box 0 0 52 52
use contact_32  contact_32_23
timestamp 1574592813
transform 1 0 31734 0 1 16236
box 0 0 52 52
use contact_32  contact_32_24
timestamp 1574592813
transform 1 0 31734 0 1 17138
box 0 0 52 52
use contact_32  contact_32_25
timestamp 1574592813
transform 1 0 32636 0 1 4510
box 0 0 52 52
use contact_32  contact_32_26
timestamp 1574592813
transform 1 0 31488 0 1 6970
box 0 0 52 52
use contact_32  contact_32_27
timestamp 1574592813
transform 1 0 31488 0 1 6068
box 0 0 52 52
use contact_32  contact_32_28
timestamp 1574592813
transform 1 0 30258 0 1 2050
box 0 0 52 52
use contact_32  contact_32_29
timestamp 1574592813
transform 1 0 30258 0 1 2706
box 0 0 52 52
use contact_32  contact_32_30
timestamp 1574592813
transform 1 0 28126 0 1 328
box 0 0 52 52
use contact_32  contact_32_31
timestamp 1574592813
transform 1 0 28126 0 1 1968
box 0 0 52 52
use contact_32  contact_32_32
timestamp 1574592813
transform 1 0 29766 0 1 2706
box 0 0 52 52
use contact_32  contact_32_33
timestamp 1574592813
transform 1 0 29766 0 1 2050
box 0 0 52 52
use contact_32  contact_32_34
timestamp 1574592813
transform 1 0 28126 0 1 2050
box 0 0 52 52
use contact_32  contact_32_35
timestamp 1574592813
transform 1 0 28126 0 1 2706
box 0 0 52 52
use contact_32  contact_32_36
timestamp 1574592813
transform 1 0 25994 0 1 328
box 0 0 52 52
use contact_32  contact_32_37
timestamp 1574592813
transform 1 0 25994 0 1 1968
box 0 0 52 52
use contact_32  contact_32_38
timestamp 1574592813
transform 1 0 26076 0 1 2050
box 0 0 52 52
use contact_32  contact_32_39
timestamp 1574592813
transform 1 0 26076 0 1 2706
box 0 0 52 52
use contact_32  contact_32_40
timestamp 1574592813
transform 1 0 24026 0 1 2050
box 0 0 52 52
use contact_32  contact_32_41
timestamp 1574592813
transform 1 0 24026 0 1 2706
box 0 0 52 52
use contact_32  contact_32_42
timestamp 1574592813
transform 1 0 22058 0 1 328
box 0 0 52 52
use contact_32  contact_32_43
timestamp 1574592813
transform 1 0 22058 0 1 984
box 0 0 52 52
use contact_32  contact_32_44
timestamp 1574592813
transform 1 0 23534 0 1 2706
box 0 0 52 52
use contact_32  contact_32_45
timestamp 1574592813
transform 1 0 23534 0 1 2050
box 0 0 52 52
use contact_32  contact_32_46
timestamp 1574592813
transform 1 0 21976 0 1 1066
box 0 0 52 52
use contact_32  contact_32_47
timestamp 1574592813
transform 1 0 21976 0 1 1968
box 0 0 52 52
use contact_32  contact_32_48
timestamp 1574592813
transform 1 0 21566 0 1 2050
box 0 0 52 52
use contact_32  contact_32_49
timestamp 1574592813
transform 1 0 21566 0 1 2706
box 0 0 52 52
use contact_32  contact_32_50
timestamp 1574592813
transform 1 0 20828 0 1 328
box 0 0 52 52
use contact_32  contact_32_51
timestamp 1574592813
transform 1 0 20828 0 1 984
box 0 0 52 52
use contact_32  contact_32_52
timestamp 1574592813
transform 1 0 19598 0 1 328
box 0 0 52 52
use contact_32  contact_32_53
timestamp 1574592813
transform 1 0 19598 0 1 984
box 0 0 52 52
use contact_32  contact_32_54
timestamp 1574592813
transform 1 0 19844 0 1 1968
box 0 0 52 52
use contact_32  contact_32_55
timestamp 1574592813
transform 1 0 19844 0 1 1066
box 0 0 52 52
use contact_32  contact_32_56
timestamp 1574592813
transform 1 0 19844 0 1 2050
box 0 0 52 52
use contact_32  contact_32_57
timestamp 1574592813
transform 1 0 19844 0 1 2706
box 0 0 52 52
use contact_32  contact_32_58
timestamp 1574592813
transform 1 0 18614 0 1 328
box 0 0 52 52
use contact_32  contact_32_59
timestamp 1574592813
transform 1 0 18614 0 1 984
box 0 0 52 52
use contact_32  contact_32_60
timestamp 1574592813
transform 1 0 17630 0 1 328
box 0 0 52 52
use contact_32  contact_32_61
timestamp 1574592813
transform 1 0 17630 0 1 984
box 0 0 52 52
use contact_32  contact_32_62
timestamp 1574592813
transform 1 0 17630 0 1 1968
box 0 0 52 52
use contact_32  contact_32_63
timestamp 1574592813
transform 1 0 17630 0 1 1066
box 0 0 52 52
use contact_32  contact_32_64
timestamp 1574592813
transform 1 0 17794 0 1 2050
box 0 0 52 52
use contact_32  contact_32_65
timestamp 1574592813
transform 1 0 17794 0 1 2706
box 0 0 52 52
use contact_32  contact_32_66
timestamp 1574592813
transform 1 0 16318 0 1 328
box 0 0 52 52
use contact_32  contact_32_67
timestamp 1574592813
transform 1 0 16318 0 1 984
box 0 0 52 52
use contact_32  contact_32_68
timestamp 1574592813
transform 1 0 15498 0 1 2050
box 0 0 52 52
use contact_32  contact_32_69
timestamp 1574592813
transform 1 0 15498 0 1 2706
box 0 0 52 52
use contact_32  contact_32_70
timestamp 1574592813
transform 1 0 15088 0 1 328
box 0 0 52 52
use contact_32  contact_32_71
timestamp 1574592813
transform 1 0 15088 0 1 984
box 0 0 52 52
use contact_32  contact_32_72
timestamp 1574592813
transform 1 0 15662 0 1 1968
box 0 0 52 52
use contact_32  contact_32_73
timestamp 1574592813
transform 1 0 15662 0 1 1066
box 0 0 52 52
use contact_32  contact_32_74
timestamp 1574592813
transform 1 0 14596 0 1 13202
box 0 0 52 52
use contact_32  contact_32_75
timestamp 1574592813
transform 1 0 14596 0 1 14104
box 0 0 52 52
use contact_32  contact_32_76
timestamp 1574592813
transform 1 0 14514 0 1 18286
box 0 0 52 52
use contact_32  contact_32_77
timestamp 1574592813
transform 1 0 14514 0 1 19188
box 0 0 52 52
use contact_32  contact_32_78
timestamp 1574592813
transform 1 0 14514 0 1 23288
box 0 0 52 52
use contact_32  contact_32_79
timestamp 1574592813
transform 1 0 14514 0 1 22304
box 0 0 52 52
use contact_32  contact_32_80
timestamp 1574592813
transform 1 0 14514 0 1 11152
box 0 0 52 52
use contact_32  contact_32_81
timestamp 1574592813
transform 1 0 14514 0 1 12054
box 0 0 52 52
use contact_32  contact_32_82
timestamp 1574592813
transform 1 0 13858 0 1 9020
box 0 0 52 52
use contact_32  contact_32_83
timestamp 1574592813
transform 1 0 13858 0 1 8118
box 0 0 52 52
use contact_32  contact_32_84
timestamp 1574592813
transform 1 0 13940 0 1 19270
box 0 0 52 52
use contact_32  contact_32_85
timestamp 1574592813
transform 1 0 13940 0 1 20254
box 0 0 52 52
use contact_32  contact_32_86
timestamp 1574592813
transform 1 0 14022 0 1 17138
box 0 0 52 52
use contact_32  contact_32_87
timestamp 1574592813
transform 1 0 14022 0 1 16236
box 0 0 52 52
use contact_32  contact_32_88
timestamp 1574592813
transform 1 0 14268 0 1 6150
box 0 0 52 52
use contact_32  contact_32_89
timestamp 1574592813
transform 1 0 14268 0 1 6970
box 0 0 52 52
use contact_32  contact_32_90
timestamp 1574592813
transform 1 0 13940 0 1 8036
box 0 0 52 52
use contact_32  contact_32_91
timestamp 1574592813
transform 1 0 13940 0 1 7052
box 0 0 52 52
use contact_32  contact_32_92
timestamp 1574592813
transform 1 0 14022 0 1 16154
box 0 0 52 52
use contact_32  contact_32_93
timestamp 1574592813
transform 1 0 14022 0 1 15252
box 0 0 52 52
use contact_32  contact_32_94
timestamp 1574592813
transform 1 0 14022 0 1 15170
box 0 0 52 52
use contact_32  contact_32_95
timestamp 1574592813
transform 1 0 14022 0 1 14186
box 0 0 52 52
use contact_32  contact_32_96
timestamp 1574592813
transform 1 0 14104 0 1 17220
box 0 0 52 52
use contact_32  contact_32_97
timestamp 1574592813
transform 1 0 14104 0 1 18204
box 0 0 52 52
use contact_32  contact_32_98
timestamp 1574592813
transform 1 0 13858 0 1 20336
box 0 0 52 52
use contact_32  contact_32_99
timestamp 1574592813
transform 1 0 13858 0 1 21238
box 0 0 52 52
use contact_32  contact_32_100
timestamp 1574592813
transform 1 0 14022 0 1 22222
box 0 0 52 52
use contact_32  contact_32_101
timestamp 1574592813
transform 1 0 14022 0 1 21320
box 0 0 52 52
use contact_32  contact_32_102
timestamp 1574592813
transform 1 0 14022 0 1 11070
box 0 0 52 52
use contact_32  contact_32_103
timestamp 1574592813
transform 1 0 14022 0 1 10168
box 0 0 52 52
use contact_32  contact_32_104
timestamp 1574592813
transform 1 0 14022 0 1 13120
box 0 0 52 52
use contact_32  contact_32_105
timestamp 1574592813
transform 1 0 14022 0 1 12136
box 0 0 52 52
use contact_32  contact_32_106
timestamp 1574592813
transform 1 0 13940 0 1 328
box 0 0 52 52
use contact_32  contact_32_107
timestamp 1574592813
transform 1 0 13940 0 1 984
box 0 0 52 52
use contact_32  contact_32_108
timestamp 1574592813
transform 1 0 12792 0 1 328
box 0 0 52 52
use contact_32  contact_32_109
timestamp 1574592813
transform 1 0 12792 0 1 984
box 0 0 52 52
use contact_32  contact_32_110
timestamp 1574592813
transform 1 0 12792 0 1 21238
box 0 0 52 52
use contact_32  contact_32_111
timestamp 1574592813
transform 1 0 12792 0 1 20336
box 0 0 52 52
use contact_32  contact_32_112
timestamp 1574592813
transform 1 0 12628 0 1 11152
box 0 0 52 52
use contact_32  contact_32_113
timestamp 1574592813
transform 1 0 12628 0 1 12054
box 0 0 52 52
use contact_32  contact_32_114
timestamp 1574592813
transform 1 0 12874 0 1 12136
box 0 0 52 52
use contact_32  contact_32_115
timestamp 1574592813
transform 1 0 12874 0 1 13120
box 0 0 52 52
use contact_32  contact_32_116
timestamp 1574592813
transform 1 0 12628 0 1 7052
box 0 0 52 52
use contact_32  contact_32_117
timestamp 1574592813
transform 1 0 12628 0 1 8036
box 0 0 52 52
use contact_32  contact_32_118
timestamp 1574592813
transform 1 0 12628 0 1 9020
box 0 0 52 52
use contact_32  contact_32_119
timestamp 1574592813
transform 1 0 12628 0 1 8118
box 0 0 52 52
use contact_32  contact_32_120
timestamp 1574592813
transform 1 0 12792 0 1 21320
box 0 0 52 52
use contact_32  contact_32_121
timestamp 1574592813
transform 1 0 12792 0 1 22222
box 0 0 52 52
use contact_32  contact_32_122
timestamp 1574592813
transform 1 0 12792 0 1 13202
box 0 0 52 52
use contact_32  contact_32_123
timestamp 1574592813
transform 1 0 12792 0 1 14104
box 0 0 52 52
use contact_32  contact_32_124
timestamp 1574592813
transform 1 0 12792 0 1 15170
box 0 0 52 52
use contact_32  contact_32_125
timestamp 1574592813
transform 1 0 12792 0 1 14186
box 0 0 52 52
use contact_32  contact_32_126
timestamp 1574592813
transform 1 0 12874 0 1 15252
box 0 0 52 52
use contact_32  contact_32_127
timestamp 1574592813
transform 1 0 12874 0 1 16154
box 0 0 52 52
use contact_32  contact_32_128
timestamp 1574592813
transform 1 0 12792 0 1 11070
box 0 0 52 52
use contact_32  contact_32_129
timestamp 1574592813
transform 1 0 12792 0 1 10168
box 0 0 52 52
use contact_32  contact_32_130
timestamp 1574592813
transform 1 0 12628 0 1 9102
box 0 0 52 52
use contact_32  contact_32_131
timestamp 1574592813
transform 1 0 12628 0 1 10086
box 0 0 52 52
use contact_32  contact_32_132
timestamp 1574592813
transform 1 0 12792 0 1 18286
box 0 0 52 52
use contact_32  contact_32_133
timestamp 1574592813
transform 1 0 12792 0 1 19188
box 0 0 52 52
use contact_32  contact_32_134
timestamp 1574592813
transform 1 0 12792 0 1 20254
box 0 0 52 52
use contact_32  contact_32_135
timestamp 1574592813
transform 1 0 12792 0 1 19270
box 0 0 52 52
use contact_32  contact_32_136
timestamp 1574592813
transform 1 0 12792 0 1 18204
box 0 0 52 52
use contact_32  contact_32_137
timestamp 1574592813
transform 1 0 12792 0 1 17220
box 0 0 52 52
use contact_32  contact_32_138
timestamp 1574592813
transform 1 0 12628 0 1 16236
box 0 0 52 52
use contact_32  contact_32_139
timestamp 1574592813
transform 1 0 12628 0 1 17138
box 0 0 52 52
use contact_32  contact_32_140
timestamp 1574592813
transform 1 0 12710 0 1 24518
box 0 0 52 52
use contact_32  contact_32_141
timestamp 1574592813
transform 1 0 12710 0 1 23370
box 0 0 52 52
use contact_32  contact_32_142
timestamp 1574592813
transform 1 0 12792 0 1 22304
box 0 0 52 52
use contact_32  contact_32_143
timestamp 1574592813
transform 1 0 12792 0 1 23288
box 0 0 52 52
use contact_32  contact_32_144
timestamp 1574592813
transform 1 0 11644 0 1 328
box 0 0 52 52
use contact_32  contact_32_145
timestamp 1574592813
transform 1 0 11644 0 1 984
box 0 0 52 52
use contact_32  contact_32_146
timestamp 1574592813
transform 1 0 11398 0 1 3034
box 0 0 52 52
use contact_32  contact_32_147
timestamp 1574592813
transform 1 0 11398 0 1 2296
box 0 0 52 52
use contact_32  contact_32_148
timestamp 1574592813
transform 1 0 11398 0 1 5494
box 0 0 52 52
use contact_32  contact_32_149
timestamp 1574592813
transform 1 0 11398 0 1 4756
box 0 0 52 52
use contact_32  contact_32_150
timestamp 1574592813
transform 1 0 11398 0 1 3116
box 0 0 52 52
use contact_32  contact_32_151
timestamp 1574592813
transform 1 0 11398 0 1 3854
box 0 0 52 52
use contact_32  contact_32_152
timestamp 1574592813
transform 1 0 11398 0 1 4674
box 0 0 52 52
use contact_32  contact_32_153
timestamp 1574592813
transform 1 0 11398 0 1 3936
box 0 0 52 52
use contact_32  contact_32_154
timestamp 1574592813
transform 1 0 10496 0 1 328
box 0 0 52 52
use contact_32  contact_32_155
timestamp 1574592813
transform 1 0 10496 0 1 984
box 0 0 52 52
use contact_32  contact_32_156
timestamp 1574592813
transform 1 0 10414 0 1 9102
box 0 0 52 52
use contact_32  contact_32_157
timestamp 1574592813
transform 1 0 10414 0 1 10086
box 0 0 52 52
use contact_32  contact_32_158
timestamp 1574592813
transform 1 0 10414 0 1 12136
box 0 0 52 52
use contact_32  contact_32_159
timestamp 1574592813
transform 1 0 10414 0 1 13120
box 0 0 52 52
use contact_32  contact_32_160
timestamp 1574592813
transform 1 0 10496 0 1 3854
box 0 0 52 52
use contact_32  contact_32_161
timestamp 1574592813
transform 1 0 10496 0 1 3116
box 0 0 52 52
use contact_32  contact_32_162
timestamp 1574592813
transform 1 0 10250 0 1 5494
box 0 0 52 52
use contact_32  contact_32_163
timestamp 1574592813
transform 1 0 10250 0 1 4756
box 0 0 52 52
use contact_32  contact_32_164
timestamp 1574592813
transform 1 0 10332 0 1 3936
box 0 0 52 52
use contact_32  contact_32_165
timestamp 1574592813
transform 1 0 10332 0 1 4674
box 0 0 52 52
use contact_32  contact_32_166
timestamp 1574592813
transform 1 0 10496 0 1 1066
box 0 0 52 52
use contact_32  contact_32_167
timestamp 1574592813
transform 1 0 10496 0 1 2214
box 0 0 52 52
use contact_32  contact_32_168
timestamp 1574592813
transform 1 0 10250 0 1 3034
box 0 0 52 52
use contact_32  contact_32_169
timestamp 1574592813
transform 1 0 10250 0 1 2296
box 0 0 52 52
use contact_32  contact_32_170
timestamp 1574592813
transform 1 0 10250 0 1 5576
box 0 0 52 52
use contact_32  contact_32_171
timestamp 1574592813
transform 1 0 10250 0 1 6970
box 0 0 52 52
use contact_32  contact_32_172
timestamp 1574592813
transform 1 0 9840 0 1 7052
box 0 0 52 52
use contact_32  contact_32_173
timestamp 1574592813
transform 1 0 9840 0 1 8036
box 0 0 52 52
use contact_32  contact_32_174
timestamp 1574592813
transform 1 0 9840 0 1 8118
box 0 0 52 52
use contact_32  contact_32_175
timestamp 1574592813
transform 1 0 9840 0 1 9020
box 0 0 52 52
use contact_32  contact_32_176
timestamp 1574592813
transform 1 0 9594 0 1 14104
box 0 0 52 52
use contact_32  contact_32_177
timestamp 1574592813
transform 1 0 9594 0 1 13202
box 0 0 52 52
use contact_32  contact_32_178
timestamp 1574592813
transform 1 0 9512 0 1 11152
box 0 0 52 52
use contact_32  contact_32_179
timestamp 1574592813
transform 1 0 9512 0 1 12054
box 0 0 52 52
use contact_32  contact_32_180
timestamp 1574592813
transform 1 0 9512 0 1 11070
box 0 0 52 52
use contact_32  contact_32_181
timestamp 1574592813
transform 1 0 9512 0 1 10168
box 0 0 52 52
use contact_32  contact_32_182
timestamp 1574592813
transform 1 0 8118 0 1 14186
box 0 0 52 52
use contact_32  contact_32_183
timestamp 1574592813
transform 1 0 8118 0 1 14924
box 0 0 52 52
use contact_32  contact_32_184
timestamp 1574592813
transform 1 0 7954 0 1 15744
box 0 0 52 52
use contact_32  contact_32_185
timestamp 1574592813
transform 1 0 7954 0 1 15006
box 0 0 52 52
use contact_32  contact_32_186
timestamp 1574592813
transform 1 0 2460 0 1 6396
box 0 0 52 52
use contact_32  contact_32_187
timestamp 1574592813
transform 1 0 2460 0 1 7134
box 0 0 52 52
use contact_32  contact_32_188
timestamp 1574592813
transform 1 0 328 0 1 7216
box 0 0 52 52
use contact_32  contact_32_189
timestamp 1574592813
transform 1 0 1640 0 1 7954
box 0 0 52 52
use contact_32  contact_32_190
timestamp 1574592813
transform 1 0 1640 0 1 7216
box 0 0 52 52
use contact_32  contact_32_191
timestamp 1574592813
transform 1 0 1804 0 1 4756
box 0 0 52 52
use contact_32  contact_32_192
timestamp 1574592813
transform 1 0 1804 0 1 5494
box 0 0 52 52
use contact_32  contact_32_193
timestamp 1574592813
transform 1 0 1722 0 1 6314
box 0 0 52 52
use contact_32  contact_32_194
timestamp 1574592813
transform 1 0 1722 0 1 5576
box 0 0 52 52
use contact_32  contact_32_195
timestamp 1574592813
transform 1 0 328 0 1 3444
box 0 0 52 52
use contact_32  contact_32_196
timestamp 1574592813
transform 1 0 1066 0 1 3444
box 0 0 52 52
use contact_32  contact_32_197
timestamp 1574592813
transform 1 0 1066 0 1 2706
box 0 0 52 52
use contact_32  contact_32_198
timestamp 1574592813
transform 1 0 32226 0 1 19762
box 0 0 52 52
use contact_32  contact_32_199
timestamp 1574592813
transform 1 0 32226 0 1 17794
box 0 0 52 52
use contact_32  contact_32_200
timestamp 1574592813
transform 1 0 32226 0 1 8528
box 0 0 52 52
use contact_32  contact_32_201
timestamp 1574592813
transform 1 0 32226 0 1 15662
box 0 0 52 52
use contact_32  contact_32_202
timestamp 1574592813
transform 1 0 32226 0 1 6478
box 0 0 52 52
use contact_32  contact_32_203
timestamp 1574592813
transform 1 0 32226 0 1 21812
box 0 0 52 52
use contact_32  contact_32_204
timestamp 1574592813
transform 1 0 32226 0 1 20746
box 0 0 52 52
use contact_32  contact_32_205
timestamp 1574592813
transform 1 0 32226 0 1 14678
box 0 0 52 52
use contact_32  contact_32_206
timestamp 1574592813
transform 1 0 32226 0 1 13612
box 0 0 52 52
use contact_32  contact_32_207
timestamp 1574592813
transform 1 0 32226 0 1 12710
box 0 0 52 52
use contact_32  contact_32_208
timestamp 1574592813
transform 1 0 32226 0 1 22796
box 0 0 52 52
use contact_32  contact_32_209
timestamp 1574592813
transform 1 0 32226 0 1 9594
box 0 0 52 52
use contact_32  contact_32_210
timestamp 1574592813
transform 1 0 32226 0 1 10660
box 0 0 52 52
use contact_32  contact_32_211
timestamp 1574592813
transform 1 0 32226 0 1 18696
box 0 0 52 52
use contact_32  contact_32_212
timestamp 1574592813
transform 1 0 32226 0 1 7544
box 0 0 52 52
use contact_32  contact_32_213
timestamp 1574592813
transform 1 0 32226 0 1 16728
box 0 0 52 52
use contact_32  contact_32_214
timestamp 1574592813
transform 1 0 32226 0 1 11562
box 0 0 52 52
use contact_32  contact_32_215
timestamp 1574592813
transform 1 0 31160 0 1 24108
box 0 0 52 52
use contact_32  contact_32_216
timestamp 1574592813
transform 1 0 31160 0 1 23862
box 0 0 52 52
use contact_32  contact_32_217
timestamp 1574592813
transform 1 0 30176 0 1 2624
box 0 0 52 52
use contact_32  contact_32_218
timestamp 1574592813
transform 1 0 30176 0 1 3198
box 0 0 52 52
use contact_32  contact_32_219
timestamp 1574592813
transform 1 0 29684 0 1 3198
box 0 0 52 52
use contact_32  contact_32_220
timestamp 1574592813
transform 1 0 29684 0 1 2624
box 0 0 52 52
use contact_32  contact_32_221
timestamp 1574592813
transform 1 0 28044 0 1 2624
box 0 0 52 52
use contact_32  contact_32_222
timestamp 1574592813
transform 1 0 28044 0 1 3198
box 0 0 52 52
use contact_32  contact_32_223
timestamp 1574592813
transform 1 0 27634 0 1 3198
box 0 0 52 52
use contact_32  contact_32_224
timestamp 1574592813
transform 1 0 27634 0 1 2624
box 0 0 52 52
use contact_32  contact_32_225
timestamp 1574592813
transform 1 0 25994 0 1 2624
box 0 0 52 52
use contact_32  contact_32_226
timestamp 1574592813
transform 1 0 25994 0 1 3198
box 0 0 52 52
use contact_32  contact_32_227
timestamp 1574592813
transform 1 0 25174 0 1 24108
box 0 0 52 52
use contact_32  contact_32_228
timestamp 1574592813
transform 1 0 25174 0 1 23862
box 0 0 52 52
use contact_32  contact_32_229
timestamp 1574592813
transform 1 0 25584 0 1 3198
box 0 0 52 52
use contact_32  contact_32_230
timestamp 1574592813
transform 1 0 25584 0 1 2624
box 0 0 52 52
use contact_32  contact_32_231
timestamp 1574592813
transform 1 0 23944 0 1 24108
box 0 0 52 52
use contact_32  contact_32_232
timestamp 1574592813
transform 1 0 23944 0 1 23862
box 0 0 52 52
use contact_32  contact_32_233
timestamp 1574592813
transform 1 0 23944 0 1 2624
box 0 0 52 52
use contact_32  contact_32_234
timestamp 1574592813
transform 1 0 23944 0 1 3198
box 0 0 52 52
use contact_32  contact_32_235
timestamp 1574592813
transform 1 0 22878 0 1 24108
box 0 0 52 52
use contact_32  contact_32_236
timestamp 1574592813
transform 1 0 22878 0 1 23862
box 0 0 52 52
use contact_32  contact_32_237
timestamp 1574592813
transform 1 0 22140 0 1 738
box 0 0 52 52
use contact_32  contact_32_238
timestamp 1574592813
transform 1 0 22140 0 1 1312
box 0 0 52 52
use contact_32  contact_32_239
timestamp 1574592813
transform 1 0 23452 0 1 3198
box 0 0 52 52
use contact_32  contact_32_240
timestamp 1574592813
transform 1 0 23452 0 1 2624
box 0 0 52 52
use contact_32  contact_32_241
timestamp 1574592813
transform 1 0 22058 0 1 1476
box 0 0 52 52
use contact_32  contact_32_242
timestamp 1574592813
transform 1 0 22058 0 1 2542
box 0 0 52 52
use contact_32  contact_32_243
timestamp 1574592813
transform 1 0 21894 0 1 2624
box 0 0 52 52
use contact_32  contact_32_244
timestamp 1574592813
transform 1 0 21894 0 1 3198
box 0 0 52 52
use contact_32  contact_32_245
timestamp 1574592813
transform 1 0 20910 0 1 738
box 0 0 52 52
use contact_32  contact_32_246
timestamp 1574592813
transform 1 0 20910 0 1 1312
box 0 0 52 52
use contact_32  contact_32_247
timestamp 1574592813
transform 1 0 20500 0 1 24108
box 0 0 52 52
use contact_32  contact_32_248
timestamp 1574592813
transform 1 0 20500 0 1 23862
box 0 0 52 52
use contact_32  contact_32_249
timestamp 1574592813
transform 1 0 19762 0 1 738
box 0 0 52 52
use contact_32  contact_32_250
timestamp 1574592813
transform 1 0 19762 0 1 1312
box 0 0 52 52
use contact_32  contact_32_251
timestamp 1574592813
transform 1 0 19762 0 1 2542
box 0 0 52 52
use contact_32  contact_32_252
timestamp 1574592813
transform 1 0 19762 0 1 1476
box 0 0 52 52
use contact_32  contact_32_253
timestamp 1574592813
transform 1 0 19762 0 1 2624
box 0 0 52 52
use contact_32  contact_32_254
timestamp 1574592813
transform 1 0 19762 0 1 3198
box 0 0 52 52
use contact_32  contact_32_255
timestamp 1574592813
transform 1 0 18532 0 1 738
box 0 0 52 52
use contact_32  contact_32_256
timestamp 1574592813
transform 1 0 18532 0 1 1312
box 0 0 52 52
use contact_32  contact_32_257
timestamp 1574592813
transform 1 0 17302 0 1 738
box 0 0 52 52
use contact_32  contact_32_258
timestamp 1574592813
transform 1 0 17302 0 1 1312
box 0 0 52 52
use contact_32  contact_32_259
timestamp 1574592813
transform 1 0 17712 0 1 2542
box 0 0 52 52
use contact_32  contact_32_260
timestamp 1574592813
transform 1 0 17712 0 1 1476
box 0 0 52 52
use contact_32  contact_32_261
timestamp 1574592813
transform 1 0 17712 0 1 2624
box 0 0 52 52
use contact_32  contact_32_262
timestamp 1574592813
transform 1 0 17712 0 1 3198
box 0 0 52 52
use contact_32  contact_32_263
timestamp 1574592813
transform 1 0 16236 0 1 738
box 0 0 52 52
use contact_32  contact_32_264
timestamp 1574592813
transform 1 0 16236 0 1 1312
box 0 0 52 52
use contact_32  contact_32_265
timestamp 1574592813
transform 1 0 16072 0 1 24108
box 0 0 52 52
use contact_32  contact_32_266
timestamp 1574592813
transform 1 0 16072 0 1 23862
box 0 0 52 52
use contact_32  contact_32_267
timestamp 1574592813
transform 1 0 16236 0 1 1476
box 0 0 52 52
use contact_32  contact_32_268
timestamp 1574592813
transform 1 0 16236 0 1 2542
box 0 0 52 52
use contact_32  contact_32_269
timestamp 1574592813
transform 1 0 15662 0 1 2624
box 0 0 52 52
use contact_32  contact_32_270
timestamp 1574592813
transform 1 0 15662 0 1 3198
box 0 0 52 52
use contact_32  contact_32_271
timestamp 1574592813
transform 1 0 15006 0 1 738
box 0 0 52 52
use contact_32  contact_32_272
timestamp 1574592813
transform 1 0 15006 0 1 1312
box 0 0 52 52
use contact_32  contact_32_273
timestamp 1574592813
transform 1 0 14514 0 1 24108
box 0 0 52 52
use contact_32  contact_32_274
timestamp 1574592813
transform 1 0 14514 0 1 23862
box 0 0 52 52
use contact_32  contact_32_275
timestamp 1574592813
transform 1 0 14514 0 1 13612
box 0 0 52 52
use contact_32  contact_32_276
timestamp 1574592813
transform 1 0 14514 0 1 12710
box 0 0 52 52
use contact_32  contact_32_277
timestamp 1574592813
transform 1 0 14596 0 1 14678
box 0 0 52 52
use contact_32  contact_32_278
timestamp 1574592813
transform 1 0 14596 0 1 15662
box 0 0 52 52
use contact_32  contact_32_279
timestamp 1574592813
transform 1 0 14678 0 1 5822
box 0 0 52 52
use contact_32  contact_32_280
timestamp 1574592813
transform 1 0 14678 0 1 6478
box 0 0 52 52
use contact_32  contact_32_281
timestamp 1574592813
transform 1 0 14596 0 1 19680
box 0 0 52 52
use contact_32  contact_32_282
timestamp 1574592813
transform 1 0 14596 0 1 18778
box 0 0 52 52
use contact_32  contact_32_283
timestamp 1574592813
transform 1 0 14596 0 1 6560
box 0 0 52 52
use contact_32  contact_32_284
timestamp 1574592813
transform 1 0 14596 0 1 7462
box 0 0 52 52
use contact_32  contact_32_285
timestamp 1574592813
transform 1 0 13940 0 1 16646
box 0 0 52 52
use contact_32  contact_32_286
timestamp 1574592813
transform 1 0 13940 0 1 15744
box 0 0 52 52
use contact_32  contact_32_287
timestamp 1574592813
transform 1 0 13940 0 1 16728
box 0 0 52 52
use contact_32  contact_32_288
timestamp 1574592813
transform 1 0 13940 0 1 17712
box 0 0 52 52
use contact_32  contact_32_289
timestamp 1574592813
transform 1 0 14022 0 1 17794
box 0 0 52 52
use contact_32  contact_32_290
timestamp 1574592813
transform 1 0 14022 0 1 18696
box 0 0 52 52
use contact_32  contact_32_291
timestamp 1574592813
transform 1 0 14022 0 1 23780
box 0 0 52 52
use contact_32  contact_32_292
timestamp 1574592813
transform 1 0 14022 0 1 22878
box 0 0 52 52
use contact_32  contact_32_293
timestamp 1574592813
transform 1 0 13940 0 1 21730
box 0 0 52 52
use contact_32  contact_32_294
timestamp 1574592813
transform 1 0 13940 0 1 20828
box 0 0 52 52
use contact_32  contact_32_295
timestamp 1574592813
transform 1 0 14022 0 1 19762
box 0 0 52 52
use contact_32  contact_32_296
timestamp 1574592813
transform 1 0 14022 0 1 20746
box 0 0 52 52
use contact_32  contact_32_297
timestamp 1574592813
transform 1 0 13940 0 1 9512
box 0 0 52 52
use contact_32  contact_32_298
timestamp 1574592813
transform 1 0 13940 0 1 8610
box 0 0 52 52
use contact_32  contact_32_299
timestamp 1574592813
transform 1 0 14022 0 1 7544
box 0 0 52 52
use contact_32  contact_32_300
timestamp 1574592813
transform 1 0 14022 0 1 8528
box 0 0 52 52
use contact_32  contact_32_301
timestamp 1574592813
transform 1 0 13940 0 1 14596
box 0 0 52 52
use contact_32  contact_32_302
timestamp 1574592813
transform 1 0 13940 0 1 13694
box 0 0 52 52
use contact_32  contact_32_303
timestamp 1574592813
transform 1 0 13940 0 1 9594
box 0 0 52 52
use contact_32  contact_32_304
timestamp 1574592813
transform 1 0 13940 0 1 10578
box 0 0 52 52
use contact_32  contact_32_305
timestamp 1574592813
transform 1 0 13940 0 1 11562
box 0 0 52 52
use contact_32  contact_32_306
timestamp 1574592813
transform 1 0 13940 0 1 10660
box 0 0 52 52
use contact_32  contact_32_307
timestamp 1574592813
transform 1 0 13940 0 1 11644
box 0 0 52 52
use contact_32  contact_32_308
timestamp 1574592813
transform 1 0 13940 0 1 12628
box 0 0 52 52
use contact_32  contact_32_309
timestamp 1574592813
transform 1 0 13858 0 1 738
box 0 0 52 52
use contact_32  contact_32_310
timestamp 1574592813
transform 1 0 13858 0 1 1312
box 0 0 52 52
use contact_32  contact_32_311
timestamp 1574592813
transform 1 0 12710 0 1 738
box 0 0 52 52
use contact_32  contact_32_312
timestamp 1574592813
transform 1 0 12710 0 1 1312
box 0 0 52 52
use contact_32  contact_32_313
timestamp 1574592813
transform 1 0 12792 0 1 6724
box 0 0 52 52
use contact_32  contact_32_314
timestamp 1574592813
transform 1 0 12792 0 1 7462
box 0 0 52 52
use contact_32  contact_32_315
timestamp 1574592813
transform 1 0 12710 0 1 7544
box 0 0 52 52
use contact_32  contact_32_316
timestamp 1574592813
transform 1 0 12710 0 1 8528
box 0 0 52 52
use contact_32  contact_32_317
timestamp 1574592813
transform 1 0 12710 0 1 18778
box 0 0 52 52
use contact_32  contact_32_318
timestamp 1574592813
transform 1 0 12710 0 1 19680
box 0 0 52 52
use contact_32  contact_32_319
timestamp 1574592813
transform 1 0 12710 0 1 10660
box 0 0 52 52
use contact_32  contact_32_320
timestamp 1574592813
transform 1 0 12710 0 1 11562
box 0 0 52 52
use contact_32  contact_32_321
timestamp 1574592813
transform 1 0 12710 0 1 13694
box 0 0 52 52
use contact_32  contact_32_322
timestamp 1574592813
transform 1 0 12710 0 1 14596
box 0 0 52 52
use contact_32  contact_32_323
timestamp 1574592813
transform 1 0 12792 0 1 8610
box 0 0 52 52
use contact_32  contact_32_324
timestamp 1574592813
transform 1 0 12792 0 1 9512
box 0 0 52 52
use contact_32  contact_32_325
timestamp 1574592813
transform 1 0 12710 0 1 10578
box 0 0 52 52
use contact_32  contact_32_326
timestamp 1574592813
transform 1 0 12710 0 1 9594
box 0 0 52 52
use contact_32  contact_32_327
timestamp 1574592813
transform 1 0 12792 0 1 16646
box 0 0 52 52
use contact_32  contact_32_328
timestamp 1574592813
transform 1 0 12792 0 1 15744
box 0 0 52 52
use contact_32  contact_32_329
timestamp 1574592813
transform 1 0 12710 0 1 14678
box 0 0 52 52
use contact_32  contact_32_330
timestamp 1574592813
transform 1 0 12710 0 1 15662
box 0 0 52 52
use contact_32  contact_32_331
timestamp 1574592813
transform 1 0 12710 0 1 18696
box 0 0 52 52
use contact_32  contact_32_332
timestamp 1574592813
transform 1 0 12710 0 1 17794
box 0 0 52 52
use contact_32  contact_32_333
timestamp 1574592813
transform 1 0 12710 0 1 16728
box 0 0 52 52
use contact_32  contact_32_334
timestamp 1574592813
transform 1 0 12710 0 1 17712
box 0 0 52 52
use contact_32  contact_32_335
timestamp 1574592813
transform 1 0 12710 0 1 21812
box 0 0 52 52
use contact_32  contact_32_336
timestamp 1574592813
transform 1 0 12710 0 1 22796
box 0 0 52 52
use contact_32  contact_32_337
timestamp 1574592813
transform 1 0 12710 0 1 19762
box 0 0 52 52
use contact_32  contact_32_338
timestamp 1574592813
transform 1 0 12710 0 1 20746
box 0 0 52 52
use contact_32  contact_32_339
timestamp 1574592813
transform 1 0 12710 0 1 21730
box 0 0 52 52
use contact_32  contact_32_340
timestamp 1574592813
transform 1 0 12710 0 1 20828
box 0 0 52 52
use contact_32  contact_32_341
timestamp 1574592813
transform 1 0 12710 0 1 13612
box 0 0 52 52
use contact_32  contact_32_342
timestamp 1574592813
transform 1 0 12710 0 1 12710
box 0 0 52 52
use contact_32  contact_32_343
timestamp 1574592813
transform 1 0 12792 0 1 11644
box 0 0 52 52
use contact_32  contact_32_344
timestamp 1574592813
transform 1 0 12792 0 1 12628
box 0 0 52 52
use contact_32  contact_32_345
timestamp 1574592813
transform 1 0 11562 0 1 738
box 0 0 52 52
use contact_32  contact_32_346
timestamp 1574592813
transform 1 0 11562 0 1 1312
box 0 0 52 52
use contact_32  contact_32_347
timestamp 1574592813
transform 1 0 11316 0 1 4346
box 0 0 52 52
use contact_32  contact_32_348
timestamp 1574592813
transform 1 0 11316 0 1 5166
box 0 0 52 52
use contact_32  contact_32_349
timestamp 1574592813
transform 1 0 11316 0 1 4264
box 0 0 52 52
use contact_32  contact_32_350
timestamp 1574592813
transform 1 0 11316 0 1 3526
box 0 0 52 52
use contact_32  contact_32_351
timestamp 1574592813
transform 1 0 11316 0 1 3444
box 0 0 52 52
use contact_32  contact_32_352
timestamp 1574592813
transform 1 0 11316 0 1 2706
box 0 0 52 52
use contact_32  contact_32_353
timestamp 1574592813
transform 1 0 10414 0 1 738
box 0 0 52 52
use contact_32  contact_32_354
timestamp 1574592813
transform 1 0 10414 0 1 1312
box 0 0 52 52
use contact_32  contact_32_355
timestamp 1574592813
transform 1 0 10332 0 1 13612
box 0 0 52 52
use contact_32  contact_32_356
timestamp 1574592813
transform 1 0 10332 0 1 12710
box 0 0 52 52
use contact_32  contact_32_357
timestamp 1574592813
transform 1 0 10414 0 1 4264
box 0 0 52 52
use contact_32  contact_32_358
timestamp 1574592813
transform 1 0 10414 0 1 3526
box 0 0 52 52
use contact_32  contact_32_359
timestamp 1574592813
transform 1 0 10414 0 1 4346
box 0 0 52 52
use contact_32  contact_32_360
timestamp 1574592813
transform 1 0 10414 0 1 5166
box 0 0 52 52
use contact_32  contact_32_361
timestamp 1574592813
transform 1 0 10414 0 1 1476
box 0 0 52 52
use contact_32  contact_32_362
timestamp 1574592813
transform 1 0 10414 0 1 2624
box 0 0 52 52
use contact_32  contact_32_363
timestamp 1574592813
transform 1 0 10332 0 1 3444
box 0 0 52 52
use contact_32  contact_32_364
timestamp 1574592813
transform 1 0 10332 0 1 2706
box 0 0 52 52
use contact_32  contact_32_365
timestamp 1574592813
transform 1 0 10332 0 1 5166
box 0 0 52 52
use contact_32  contact_32_366
timestamp 1574592813
transform 1 0 10332 0 1 7462
box 0 0 52 52
use contact_32  contact_32_367
timestamp 1574592813
transform 1 0 9758 0 1 7544
box 0 0 52 52
use contact_32  contact_32_368
timestamp 1574592813
transform 1 0 9758 0 1 8528
box 0 0 52 52
use contact_32  contact_32_369
timestamp 1574592813
transform 1 0 9758 0 1 8610
box 0 0 52 52
use contact_32  contact_32_370
timestamp 1574592813
transform 1 0 9758 0 1 10578
box 0 0 52 52
use contact_32  contact_32_371
timestamp 1574592813
transform 1 0 9594 0 1 10660
box 0 0 52 52
use contact_32  contact_32_372
timestamp 1574592813
transform 1 0 9594 0 1 11562
box 0 0 52 52
use contact_32  contact_32_373
timestamp 1574592813
transform 1 0 9594 0 1 12628
box 0 0 52 52
use contact_32  contact_32_374
timestamp 1574592813
transform 1 0 9594 0 1 11644
box 0 0 52 52
use contact_32  contact_32_375
timestamp 1574592813
transform 1 0 9512 0 1 13694
box 0 0 52 52
use contact_32  contact_32_376
timestamp 1574592813
transform 1 0 9512 0 1 14514
box 0 0 52 52
use contact_32  contact_32_377
timestamp 1574592813
transform 1 0 8036 0 1 14596
box 0 0 52 52
use contact_32  contact_32_378
timestamp 1574592813
transform 1 0 8036 0 1 15334
box 0 0 52 52
use contact_32  contact_32_379
timestamp 1574592813
transform 1 0 8118 0 1 15416
box 0 0 52 52
use contact_32  contact_32_380
timestamp 1574592813
transform 1 0 8118 0 1 16154
box 0 0 52 52
use contact_32  contact_32_381
timestamp 1574592813
transform 1 0 2296 0 1 7544
box 0 0 52 52
use contact_32  contact_32_382
timestamp 1574592813
transform 1 0 2296 0 1 6806
box 0 0 52 52
use contact_32  contact_32_383
timestamp 1574592813
transform 1 0 2378 0 1 6724
box 0 0 52 52
use contact_32  contact_32_384
timestamp 1574592813
transform 1 0 2378 0 1 5986
box 0 0 52 52
use contact_32  contact_32_385
timestamp 1574592813
transform 1 0 1640 0 1 5904
box 0 0 52 52
use contact_32  contact_32_386
timestamp 1574592813
transform 1 0 1640 0 1 5166
box 0 0 52 52
use contact_32  contact_32_387
timestamp 1574592813
transform 1 0 738 0 1 4264
box 0 0 52 52
use contact_32  contact_32_388
timestamp 1574592813
transform 1 0 1722 0 1 5166
box 0 0 52 52
use contact_32  contact_32_389
timestamp 1574592813
transform 1 0 1722 0 1 4346
box 0 0 52 52
use contact_32  contact_32_390
timestamp 1574592813
transform 1 0 738 0 1 3034
box 0 0 52 52
use contact_32  contact_32_391
timestamp 1574592813
transform 1 0 27880 0 1 2952
box 0 0 52 52
use contact_32  contact_32_392
timestamp 1574592813
transform 1 0 25912 0 1 2952
box 0 0 52 52
use contact_32  contact_32_393
timestamp 1574592813
transform 1 0 23780 0 1 2952
box 0 0 52 52
use contact_32  contact_32_394
timestamp 1574592813
transform 1 0 21730 0 1 2952
box 0 0 52 52
use contact_32  contact_32_395
timestamp 1574592813
transform 1 0 19680 0 1 2952
box 0 0 52 52
use contact_32  contact_32_396
timestamp 1574592813
transform 1 0 17466 0 1 2952
box 0 0 52 52
use contact_32  contact_32_397
timestamp 1574592813
transform 1 0 15580 0 1 2952
box 0 0 52 52
use contact_32  contact_32_398
timestamp 1574592813
transform 1 0 4182 0 1 2870
box 0 0 52 52
use contact_32  contact_32_399
timestamp 1574592813
transform 1 0 12300 0 1 1312
box 0 0 52 52
use contact_32  contact_32_400
timestamp 1574592813
transform 1 0 11152 0 1 1312
box 0 0 52 52
use contact_32  contact_32_401
timestamp 1574592813
transform 1 0 9922 0 1 1312
box 0 0 52 52
use contact_32  contact_32_402
timestamp 1574592813
transform 1 0 21566 0 1 1312
box 0 0 52 52
use contact_32  contact_32_403
timestamp 1574592813
transform 1 0 20418 0 1 1312
box 0 0 52 52
use contact_32  contact_32_404
timestamp 1574592813
transform 1 0 19270 0 1 1312
box 0 0 52 52
use contact_32  contact_32_405
timestamp 1574592813
transform 1 0 18040 0 1 1312
box 0 0 52 52
use contact_32  contact_32_406
timestamp 1574592813
transform 1 0 16974 0 1 1312
box 0 0 52 52
use contact_32  contact_32_407
timestamp 1574592813
transform 1 0 15744 0 1 1312
box 0 0 52 52
use contact_32  contact_32_408
timestamp 1574592813
transform 1 0 14596 0 1 1312
box 0 0 52 52
use contact_32  contact_32_409
timestamp 1574592813
transform 1 0 13448 0 1 1312
box 0 0 52 52
use contact_32  contact_32_410
timestamp 1574592813
transform 1 0 1175 0 1 7771
box 0 0 52 52
use contact_32  contact_32_411
timestamp 1574592813
transform 1 0 1175 0 1 5035
box 0 0 52 52
use contact_34  contact_34_0
timestamp 1574592870
transform 1 0 32636 0 1 246
box 0 0 52 52
use contact_34  contact_34_1
timestamp 1574592870
transform 1 0 246 0 1 24600
box 0 0 52 52
use contact_34  contact_34_2
timestamp 1574592870
transform 1 0 246 0 1 246
box 0 0 52 52
use contact_34  contact_34_3
timestamp 1574592870
transform 1 0 32718 0 1 24600
box 0 0 52 52
use contact_34  contact_34_4
timestamp 1574592870
transform 1 0 32718 0 1 246
box 0 0 52 52
use contact_34  contact_34_5
timestamp 1574592870
transform 1 0 164 0 1 246
box 0 0 52 52
use contact_34  contact_34_6
timestamp 1574592870
transform 1 0 32800 0 1 24600
box 0 0 52 52
use contact_34  contact_34_7
timestamp 1574592870
transform 1 0 328 0 1 24600
box 0 0 52 52
use contact_34  contact_34_8
timestamp 1574592870
transform 1 0 328 0 1 246
box 0 0 52 52
use contact_34  contact_34_9
timestamp 1574592870
transform 1 0 164 0 1 24682
box 0 0 52 52
use contact_34  contact_34_10
timestamp 1574592870
transform 1 0 164 0 1 328
box 0 0 52 52
use contact_34  contact_34_11
timestamp 1574592870
transform 1 0 32800 0 1 246
box 0 0 52 52
use contact_34  contact_34_12
timestamp 1574592870
transform 1 0 32636 0 1 24682
box 0 0 52 52
use contact_34  contact_34_13
timestamp 1574592870
transform 1 0 32636 0 1 328
box 0 0 52 52
use contact_34  contact_34_14
timestamp 1574592870
transform 1 0 32636 0 1 24518
box 0 0 52 52
use contact_34  contact_34_15
timestamp 1574592870
transform 1 0 246 0 1 24682
box 0 0 52 52
use contact_34  contact_34_16
timestamp 1574592870
transform 1 0 246 0 1 328
box 0 0 52 52
use contact_34  contact_34_17
timestamp 1574592870
transform 1 0 32718 0 1 24682
box 0 0 52 52
use contact_34  contact_34_18
timestamp 1574592870
transform 1 0 246 0 1 24518
box 0 0 52 52
use contact_34  contact_34_19
timestamp 1574592870
transform 1 0 246 0 1 164
box 0 0 52 52
use contact_34  contact_34_20
timestamp 1574592870
transform 1 0 32718 0 1 328
box 0 0 52 52
use contact_34  contact_34_21
timestamp 1574592870
transform 1 0 32718 0 1 24518
box 0 0 52 52
use contact_34  contact_34_22
timestamp 1574592870
transform 1 0 164 0 1 24518
box 0 0 52 52
use contact_34  contact_34_23
timestamp 1574592870
transform 1 0 32718 0 1 164
box 0 0 52 52
use contact_34  contact_34_24
timestamp 1574592870
transform 1 0 164 0 1 164
box 0 0 52 52
use contact_34  contact_34_25
timestamp 1574592870
transform 1 0 32636 0 1 164
box 0 0 52 52
use contact_34  contact_34_26
timestamp 1574592870
transform 1 0 328 0 1 24682
box 0 0 52 52
use contact_34  contact_34_27
timestamp 1574592870
transform 1 0 32800 0 1 24682
box 0 0 52 52
use contact_34  contact_34_28
timestamp 1574592870
transform 1 0 32800 0 1 328
box 0 0 52 52
use contact_34  contact_34_29
timestamp 1574592870
transform 1 0 328 0 1 328
box 0 0 52 52
use contact_34  contact_34_30
timestamp 1574592870
transform 1 0 328 0 1 24518
box 0 0 52 52
use contact_34  contact_34_31
timestamp 1574592870
transform 1 0 328 0 1 164
box 0 0 52 52
use contact_34  contact_34_32
timestamp 1574592870
transform 1 0 164 0 1 24600
box 0 0 52 52
use contact_34  contact_34_33
timestamp 1574592870
transform 1 0 32800 0 1 24518
box 0 0 52 52
use contact_34  contact_34_34
timestamp 1574592870
transform 1 0 32800 0 1 164
box 0 0 52 52
use contact_34  contact_34_35
timestamp 1574592870
transform 1 0 32636 0 1 24600
box 0 0 52 52
use contact_34  contact_34_36
timestamp 1574592870
transform 1 0 738 0 1 24190
box 0 0 52 52
use contact_34  contact_34_37
timestamp 1574592870
transform 1 0 32390 0 1 24108
box 0 0 52 52
use contact_34  contact_34_38
timestamp 1574592870
transform 1 0 738 0 1 738
box 0 0 52 52
use contact_34  contact_34_39
timestamp 1574592870
transform 1 0 32390 0 1 656
box 0 0 52 52
use contact_34  contact_34_40
timestamp 1574592870
transform 1 0 32226 0 1 24190
box 0 0 52 52
use contact_34  contact_34_41
timestamp 1574592870
transform 1 0 32308 0 1 24190
box 0 0 52 52
use contact_34  contact_34_42
timestamp 1574592870
transform 1 0 32308 0 1 738
box 0 0 52 52
use contact_34  contact_34_43
timestamp 1574592870
transform 1 0 574 0 1 738
box 0 0 52 52
use contact_34  contact_34_44
timestamp 1574592870
transform 1 0 32226 0 1 738
box 0 0 52 52
use contact_34  contact_34_45
timestamp 1574592870
transform 1 0 738 0 1 574
box 0 0 52 52
use contact_34  contact_34_46
timestamp 1574592870
transform 1 0 656 0 1 24190
box 0 0 52 52
use contact_34  contact_34_47
timestamp 1574592870
transform 1 0 32226 0 1 574
box 0 0 52 52
use contact_34  contact_34_48
timestamp 1574592870
transform 1 0 656 0 1 738
box 0 0 52 52
use contact_34  contact_34_49
timestamp 1574592870
transform 1 0 574 0 1 24190
box 0 0 52 52
use contact_34  contact_34_50
timestamp 1574592870
transform 1 0 656 0 1 574
box 0 0 52 52
use contact_34  contact_34_51
timestamp 1574592870
transform 1 0 32308 0 1 574
box 0 0 52 52
use contact_34  contact_34_52
timestamp 1574592870
transform 1 0 574 0 1 574
box 0 0 52 52
use contact_34  contact_34_53
timestamp 1574592870
transform 1 0 32390 0 1 24190
box 0 0 52 52
use contact_34  contact_34_54
timestamp 1574592870
transform 1 0 738 0 1 24272
box 0 0 52 52
use contact_34  contact_34_55
timestamp 1574592870
transform 1 0 32390 0 1 738
box 0 0 52 52
use contact_34  contact_34_56
timestamp 1574592870
transform 1 0 32390 0 1 574
box 0 0 52 52
use contact_34  contact_34_57
timestamp 1574592870
transform 1 0 656 0 1 24272
box 0 0 52 52
use contact_34  contact_34_58
timestamp 1574592870
transform 1 0 32308 0 1 24272
box 0 0 52 52
use contact_34  contact_34_59
timestamp 1574592870
transform 1 0 574 0 1 24272
box 0 0 52 52
use contact_34  contact_34_60
timestamp 1574592870
transform 1 0 738 0 1 24108
box 0 0 52 52
use contact_34  contact_34_61
timestamp 1574592870
transform 1 0 32308 0 1 24108
box 0 0 52 52
use contact_34  contact_34_62
timestamp 1574592870
transform 1 0 32308 0 1 656
box 0 0 52 52
use contact_34  contact_34_63
timestamp 1574592870
transform 1 0 32226 0 1 24272
box 0 0 52 52
use contact_34  contact_34_64
timestamp 1574592870
transform 1 0 574 0 1 24108
box 0 0 52 52
use contact_34  contact_34_65
timestamp 1574592870
transform 1 0 738 0 1 656
box 0 0 52 52
use contact_34  contact_34_66
timestamp 1574592870
transform 1 0 32226 0 1 24108
box 0 0 52 52
use contact_34  contact_34_67
timestamp 1574592870
transform 1 0 32226 0 1 656
box 0 0 52 52
use contact_34  contact_34_68
timestamp 1574592870
transform 1 0 656 0 1 24108
box 0 0 52 52
use contact_34  contact_34_69
timestamp 1574592870
transform 1 0 656 0 1 656
box 0 0 52 52
use contact_34  contact_34_70
timestamp 1574592870
transform 1 0 574 0 1 656
box 0 0 52 52
use contact_34  contact_34_71
timestamp 1574592870
transform 1 0 32390 0 1 24272
box 0 0 52 52
use control_logic_rw  control_logic_rw_0
timestamp 1574592812
transform 1 0 1146 0 1 2711
box -132 -36 7665 5304
use cr_10  cr_10_0
timestamp 1574592813
transform 1 0 8882 0 1 1912
box 1192 -673 4309 1361
use cr_11  cr_11_0
timestamp 1574592813
transform 1 0 8882 0 1 1912
box 5425 -692 20788 328
use data_dff  data_dff_0
timestamp 1574592812
transform 1 0 13410 0 1 1014
box -116 -36 9320 451
use row_addr_dff  row_addr_dff_0
timestamp 1574592812
transform 1 0 7585 0 1 14185
box -116 -36 1165 2075
<< labels >>
rlabel metal3 67 2896 67 2896 4 csb0
rlabel metal3 67 3306 67 3306 4 web0
rlabel metal4 4208 67 4208 67 4 clk0
rlabel metal4 13474 67 13474 67 4 din0[0]
rlabel metal4 14622 67 14622 67 4 din0[1]
rlabel metal4 15770 67 15770 67 4 din0[2]
rlabel metal4 17000 67 17000 67 4 din0[3]
rlabel metal4 18066 67 18066 67 4 din0[4]
rlabel metal4 19296 67 19296 67 4 din0[5]
rlabel metal4 20444 67 20444 67 4 din0[6]
rlabel metal4 21592 67 21592 67 4 din0[7]
rlabel metal4 15606 67 15606 67 4 dout0[0]
rlabel metal4 17492 67 17492 67 4 dout0[1]
rlabel metal4 19706 67 19706 67 4 dout0[2]
rlabel metal4 21756 67 21756 67 4 dout0[3]
rlabel metal4 23806 67 23806 67 4 dout0[4]
rlabel metal4 25938 67 25938 67 4 dout0[5]
rlabel metal4 27906 67 27906 67 4 dout0[6]
rlabel metal3 32949 2978 32949 2978 4 dout0[7]
rlabel metal4 9948 67 9948 67 4 addr0[0]
rlabel metal4 11178 67 11178 67 4 addr0[1]
rlabel metal4 12326 67 12326 67 4 addr0[2]
rlabel metal3 67 14458 67 14458 4 addr0[3]
rlabel metal3 67 14786 67 14786 4 addr0[4]
rlabel metal3 67 15278 67 15278 4 addr0[5]
rlabel metal3 67 15524 67 15524 4 addr0[6]
rlabel metal3 67 16016 67 16016 4 addr0[7]
rlabel metal4 32334 12449 32334 12449 4 vdd
rlabel metal3 16508 682 16508 682 4 vdd
rlabel metal3 16508 24216 16508 24216 4 vdd
rlabel metal4 682 12449 682 12449 4 vdd
rlabel metal3 16508 272 16508 272 4 gnd
rlabel metal4 32744 12449 32744 12449 4 gnd
rlabel metal4 272 12449 272 12449 4 gnd
rlabel metal3 16508 24626 16508 24626 4 gnd
<< properties >>
string FIXED_BBOX 0 0 33016 24734
<< end >>
